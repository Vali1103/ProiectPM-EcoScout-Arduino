PK   ���XR d�eu  l    cirkitFile.json��9�%�*	f������k�0���nt��.�U�g�0*ENH�(����3-�7B��e7�0U���BVJ~i~����F3'��������p�0���������7ߓ���������o���������|�~�Û��T��>�돓��n��K����׺�j&G�Q�U_�F�1irf������~���oOw��ۯ͇�?�x�q���.��4�bqҽr�v*wI�nuУ��Dw���o%���%tA �@��-��~�A�1��aR��N���sS��Н7"ta_�߈�Տ�	�������A=t�?���ݏ������U}���+ԣr)���sb58�������mx!^̆�F�������Җ��l�H!uvQ�R�.�1H-�,� �P:�t�%���0~KM�QXl���rR�xq8�G8�'��F:� �HVB���&

��((�>\l���{q��?�ݸ�DA!w�b��O$�\�r#����L6�M�X�J��@�^���B��B���DA!���&

��%6QP�,���B>`�M�KlB�Y��%6QP�,���Bw�M�Cl����N���B�;�&

���((�Sl����N���B�;�&����N���B�;�&

���((�Sl�� ����}��DA!��b��w�Mr�)6QP�}��D	�Sl����N�	]��br���Sl����N������N/��b��w.&D�ۀL��]�z��$dNF�8�D��RB�l�U���-�G4���b�~Jq��T�'*�U7�\��)O�l�x����ȸ<�ޫ<�S��I��4��>��������(|A>
��t������{3)��Q];��)�A�1u�s]:g���r���aJ*Q�l_`�4Ș�e���;&����NZ�z���]
N�)�4k���Qb�����31Оc"ؕ0���=�,=�*����������"Y�Mc�s6��O������܏�7��D��O�[j�}���I62.���8��L,�y<&���4�DY$V��,��@j�R�'󏛣T�<�Қ옔�]�r�^E��0L��1����{� ̧?X7ab�Z8�3db�Z8�3�
0Z�k���:C.
���H��BjB�qQHM���<.
����>.
��>��㢐�ͣ�<.
��<��㢐�Σ�<�]�;�*�(�� ���4r�)6�Xg&
^̶�O$��Gg\r?l��װ�=[f�svV;�5:���R2N7��̘m����l������5��*��-GEt\��d)����8usVy��&MAu�y՛�OYS�R/W��1��Ԅ�ֈ� �]gDP*��Zh/�BkV`�.O&#����+r�·F�o�u^���bf���j�q���R����[��*{"�tqO~�Dd^���y�>�LƓ��n9�Ͻuc�um���J�L2\,s��d���d��}0Z?��'�YX<I�|0Z?��v�U�ǹ����۩�>��MFU�2����#,:}��E��bJ~r��Ţr~�������H&�%�/�	�`�~0O	K{�J�����]�r���A�]�Ja�#h�E`|�W�i`�����_�r&��'�u�)���)σr��~ ��$��4ڡ�G�كPǈ��^�t��>m<��*h��jF��C��(?m<��.phF������������#,,>�`�����_-� ������u���LX|�W�Q��pЄ�G`|���8h��#0�Z��`�_-^������USH{���_-���?���ﺺ�8���#0�Z��`�ߺ�o���cM�z�뷻Ψ����{�:���+]�P ԃC,��?�t�����]�58�������~�`�����՝���C,>�{T��c%mXC���]E�z,8������ꖢ`��Q����P����,>�۸��G=X|�W7��]����n���`�_��˟�.X|�W�+�]����n���`�_�"�8��G`|usk0�qП���?8���#0���8�?p���G`|u+t0�������&�`������������,>��c����������`�������
����,>��,���X|�W� ��?����m�`���Q�V����^u҆�.p��~<!]��Ń�,>�>z��*<x�|���^A8�Y?��.p�������CV��p��G`|�x0۽=�#����r�K���S}A��su�9����G��GR�k�7�wa�ͨL��r]7�4���<��#�S�r��1���v�q�a»����o�CWhw��=8�d��)��vcy�vH��X����C��l�A;�S}6���܃���s�?�a���;��Qz��y������s�Mn7�����S#�x&,w�%��OX���;5�n��E�TX��b�}D��8�:���U.�TlY��-v��ϱ;���{V�v�"���A�F�v?6�	B��ś��A�p��D�}�8 @GS�p
O�*pD��	�� ���",�vj|�=�����_a�8���a��W؃�r��n�/�� ��,��K|�=�`���_a�8j��a��W؃�?��n�/���a�ݰ_"��Q0������G����X|7��>��8���a��W�2+�iv���!��[0�������+�A��/X|7l���Á��!Hs��臽[#��a0������_y��Pn�¡vld��<�wD|uіx�[�5"%d���m�{E~�:$ӧ)�c��aV�|Tv�y�S��=Qs�57��V��ɚ{Y��������76y����_��~�l��ꎄ�#��H(=j���#��H(?���g�~O�?#ԟ���g��3B����PV�?��?g��aPi,M�&��I;7E����»�|_�����g5�W>����Y��u�j�/{V�}��d#��Pw�>��Py�>��P{�>��P}�>��P�>����	�w0����w0����w0����w0��.�������B�Y���PV�?+ԟ��
���sB�9s�w��/��(�I��Y�d�`EЅ��	{��'�N���x�y�����L��t�\���]ҪG�h�<ы?n��u�}����-��֍!�**�SUrѩ���5�9�Q��{ݍu̼쩽��ѭ�=�G�\��"�Iz{{Yx{#�}��ۋF� ��p��l����5j�ME؍�p��7�(p�P�Q(�(�rJ9
'|Q��(�_�/
����KB�%���PI��$�_�/I���KB�e���PY��,�_�/�����B�ei�E�v��]�4񢥙-M�hi�EK�/Z�}����_�T���T���8	(��Ӏ�<�8(�JS�$��4H�l IӁ$��4!HҌ IS�$�	�4)HҬ Iӂ$��41H�� IS�$��49H�� IӃ$��4AHN�Di^��T���I�s$MБ4CG�Ist�J�R%z���ZL�Di���T�^�D/Ub�*Q��!i&�����b(��J��PH�D!i��i��QH�H!i&�����RH�L!i6�����SH�P!iF��)��TH�T!iV��i��UH�X!if�����V(_�d}m�ٞ�h��Ӕ�KΩ>u�r]�Sof�WG��|ｂ,ֽE�=$M�Pޫ��Ny����W�֩l�^�)�ݜu7��$�w�'c˽}�������Fu}o�8��	�('ɽ���?��;�C}��S4�Fn�Hud�JѤA�:LAX~h�n�'�ޢ�f��3#͝i���Θ��f��z����<��oߛ)Z��k��[�ܵ�lߛ9,�8߫�d��{�m2G5ѽ�����;��6�c���ۍ�3��uF�>'=�.�#�����X���+���we5������{3E�I͆Ꙁ�����f�X�j=�p�����6��!��{.�u�k��^���[��BH�{�Űn}�ܷ�E[NY4��c0����}�"y��� ��{'���}�<]a
��y�W� ��������H�����E��ݮ,cJ~r���H��ܫ.wVѠ�����A��DV�� ��T\�U�2�'��Ӭ��:�bYg��R����R�K��D*�:_�AZ�_�X߲p��q�u�sv���)����$;Q,��ѥa����2^�6,��GB�M��
�Txs���� X�)O�\fT���s��$�����GB���L%��e���Fuq�Jd=%?�1��+�8#Nc�u��2�΁�{n�r��-���s�z̎�l	3\	q�>��C�W&��+�����>�QX��c����x�Rpgi���s怵��5o��Y��{wgm>��6ށ���k���k̍ww��W�,�����j��e5�ό����EY��3%<	J%,���'��B|`�k/������Q�Y����|��
�|���P��h���lv7/�����n��cg�zw��u�;��{�&ޭ�2�qʼp�%��r�)�i��7����2��w�M�[�[�8gg�+���z�J�8e��3c�a���7�؛,�)��2Vd�2A�]]�^E��0���ٯ���zw���Mo9d�r�{�&c��<�6�vS��ѶK��>����G�����e��E����l7yMq��w�4"�UG%��S�%�J�40�j~r��3�j�ϼ�G��P:gWZ:��S!������������?;�������?;�;ﮀ1�F���;�^��+1G,�a+f�B�9NKn�W4���Hn��a�ӻ+q�;R��Y������X���q�E��{�繏C�S�U��8t�a95������\�rY��].s�$xp��va�Z6��w{�ŧ���U]\.c��e���y�M������|��4��j������S6�g]gba��V�Г��h�bH�H&�J���.�����ǜ�����{���SE���>���k��@�t4��B��LlM_�[.�S�#��/]~*3�~���T�<�Vs���}�a�9O�:W���<-'=��ػ"m�ۃ���/w��������p��������hDo�C�	Û��7DCz�GbhI� ѓ�8�^�Ƞٺ΍��J�������:e�p�����:�(D�(�-��q���E"�!]�D C��L0�@�����H��ƹm�%�d�@�@����aY�KV3�h�K��	4�%�zw Kz��0�|8��8ʒ^҅ L0?n`~eI/iM&�7���z�b2���Y�o��8J1���6	GY�K��	��̏�,-�£0�����q��e}�	��-̏�,�%y���6GY���s L�����q�%�������Q��r�̏[�GY�ˁ� L0?�`~eI/#�0�����q���	��Q��r�#̏;�GY�˱� L0?�`~eI/�[�0�����q�%��	J������q�%���	�����Q��rD(̏{\z��=̏�,��R��Z��	�۸XB�g������Q��/@�Zt�g/\�0?�;��u"У�CL��0�8uELD�t3-�bt��lz2���LD�C&�yN���<5�Dt^W�Dt>\2��1��LD C�uE�.©+�~���d�SW�D2Ī+�H��ƹm�%V]l�eTq1�,iN5Ȓ�Tq1�,�ꊸ�`�Q����j .&�gTq1��8��;���qF5̏���̏�,=��g���".&�GYz�+B+��".�{w0?Ψ�b��qs���Ŵ��o�RQ_ƽ�EV�g�O}�U��*g�6�"x�&�R^�X���"x5��v���+m`E0`��j���+m`E0���� +m`[���կ���5�JX�&��&zm���`����kl�_[`��R^S���JM���w�[��+5�Z�M��Q�AKm��<Nn[D2�-�A�>ж�fh-�,��6���s�P�m¯�Z5�f�ܶ	�6�BHh�Q�Ȇڠ�6hk���m"�&h�ښwn�m��ڠ�6hk���m"�&h��ZІ�6QY��m�gh�Xh�5AKm�ֺ�6ܶ�˚��6hk}In��eM�R��N��-"j��ڠ��>m�m�k��ڠ�uKm�m�5AKm����6ܶ�˚��6hkYn��eM�R��3�A뷦M\��m�m��̴�˚��6h�gm
���eM�R�u��6ܶ�˚��6h�>tm�m�5AKm�����pۨZ�Q�b��̶��l���	Zj���o؆�6qY��mݧ��m�&h�ں�dn��eM�R�u��6ܶ�˚��6h���m�m�5AKm��}L�p���eM�R�u?�6ܶ�˚��6h뾲m�m�5AKm���q�p�&_�-�A[��m�m�/�}J�&.sm�2�&.k��ڠ��.��M\�-�A[��n�m���	Zj���݆�6qY��m�ϻ�m�&h�ں/yn}���	Zj���ކ�6qY��m�'��m�&h�ں�}n��eM�R�u��6ܶ�˚��6h��m�m�5AKm��s�p��t9�&hi-��6q�o�5AKm��s-�p��t �m�m����&.�m�&h��z�HnC���	Zj����҆�6�-6AK[h!$���B����-��f�����v�f�G�4�z�ޫ��қ�zc����ބ�Xo�{�v�@���z�ޫ����z�z�Х&���z�ޫ�[�z����V��޸�q�U �-�޼�*���&�޸��=ƫ	�-�޼���V����z�ޫ��Κ�z�J�H�&�޸�=��ɸu��`�&���z�ޫ�0��ڄ\M�޾��+�"�mv���n���f�ܶ	����}��W�Er�&�j����W_a�m��	���^}�Y$�m°&ho�{�f�ܶ	Ś��}��W�Er�&k����W_a�m���	���^}�Y$�m²&ho�{�f��6A{�ޫ�3q�p�&.k����W�g���M\���{���(n�m���	���^e���d����L��9��M\v�n��0��M\���{���,��M\v�ޫ�3��p�&.k����W�g���m�[�^}�Y$�m�e��B|B������p���?N?߅d�4�Qu1�ʅ0�L>*;�<�)v]7�i��X1+b�A�x�� �!V�Jƨ$^�z	#_��0&��	#a�h�0"&��F��1*6��F��b�Q����`Tl1*��*vV�q��b�aR��N���sS������e��C����'����ĲrڛXVN;��i_bY9�J,+�=��:�x1�=����`�{>���(�|V�3������g���Y��cT|>�����|V�3�Q����g���Yo�Ũ4����F��b�Q�Ũ�bTl1*�;��F��l���j4#^T<���Qb�b�Q�è�aT�0*��GwS�$f}q{/1��x0iȳ�̣/Ns$f���������湐-0�.=<��J�,*�z�MXT'3�"3_03����3�~;�w�����/_1�8bT1*�G��#fFA�lG��#F�	��Qq¨8aT�0*N'��h���Qqƨ8cT�1*�g��3F���Qq%=PYP�C����Р̇�>4(��A��~hP�C��K��J�2y�T*��J桲y�t(�G���2zJ�(�G����zJ�(�G���2{J�(�G����{J�(�G��2|J�(�G�$��|�@z��ȁ���(�G�\��}��(�G�gҳ�٣J�@z%�ȃ��Az� =��A�?����#P����gP��@	@e 	�$P�@I@e	�$P�@�@e	�
$P.�@�@e	�$P>�@	Ae	�$PN�@IAe	�$P^���u%v=�I�$�Q#Pj�s��:�Y���_�g�%�at�f���Dv���I(?h��%�Tu�K~0Ө�^d�I	(?h@�As���������:�:?�N����7v��a���<R�
�i9��';;ESy7w�:�Q�hҠ{�0ޝ*�e�T7��i�&+=MI���SW�uyN��ma�ˁdY�3ؗKy��]MuG�Bq�c���nκ�<b9�\,+t淢M�)Vܨ�1��]gT�s�S�B1w��.���XŲrڳYVN�5��i�fY9��ݛ)�Nj6TTח~�{[z�Mc1��c����}
�j�̤�I��خ<QҪG�h�<}��{���ee��d�N���[7�ث��̢{�\t�s>�Na���Q?�ʂ�j�e��㚁h���:]�no��<��a��>N�':�²����?J`Y9}�1Ř�Ҷ��XqΨ�_������q��Db+��eey���,XV�e���pi�)��u*�~���{���*��#���:|�+�7M�<��uN)LF�h�z��=�Jz��O��i<:���XY��U���i;t�}.ZW�T��By�`�능�q���e���Ҏ��8��l�'_�������!�<��#ݗ�<����%;ڝ�K�p���<�7���Fuq�ʴlJ~�cLOz9���e�K)��M�L5��u������wS���4,G�����#[�5WFءO�M�_}��*b�����>YVN�Ʈ���U�N��_;�~(��D�L�D٥�wt�XV��MS�BC��U/՗'��YEu��m������e�����c~��F��zT�{fSf�֧�1��cY9}G,+�sL���9&ˊ;YVN�,+��z,+�kz,+�+z,+��<ՁċQ�y1)�F�祤<3������x�e#��*R��è����g���
R���/��s��� 1.fz�[��YT\��^l�2���� 3��x�R����o�;�d:�T9�ߋw�)������c	4rP��ʬ�����]�{�q��gy8V���9V�W�9V���9VNǄn����liK֫�J�2�.�j������G+��e���y�:N��p6h՗��P��<�h���yaY9�e���S^F7�!����*�MR]�V�J���p�XcY��5/�s��YV��p²��ƶ8usV�D���T�tv^�&�S�Tb���]�:�\���کn����G��)�q�Ό�b�yq��ٸ��>}OE��P"����ujs�C��网e�7��z�Vd�T��ꊶ.��d;5�`���X��K�n���)ǹ��RP��T?_���:�@)v/űr�K��h�O�b!��8�<e�Lp�u&�Ycg[����3UZFŐ\yӁT�e4��φz����VN�����:U�V��*B/���MG��9ǀe�|d��r!v�����˩����!��p͘�q��bs�rΓ��v�2b���l�]7����XXV�c��b����ݧ�������j��J���a��\�;�f�N��\�]u]m���`SWO��>N?}~�><�w�!B���B��e� ��hA2���Ȑ^""�!���B��e��dH/k�D CzY?� җ�h���ym�ۆ�m�9n�%}Yr�`��n�9o�%}I`0��7�8ʒ��)0�`>�`NeI_(L0?n`~eI_R;L��7n����Q��%�������Q��%�������Q��%������Q��%�	�a~���8ʒ������[I�-������q�%}9&�	��-̏�,��&L0?na~eI_�V�`��q��(K�r�̏;�GY*�`~eI_ζ�`��q��(K�r�̏;�GYҗ�0�`~���8ʒ��T�I������q�%}9C	�	��=̏�,���NL��&.�	����Q���+&��0?���/�ka0��x��q�%}9��	��̏3,M�Փ����X�����Rp*L)�Yk?��"�!N]�9�LD C��"&"�[;2��@�8uELD C��"&"�!N]�����d�SW�D2ĩ+b"b�q]$�k��6�o3����`��Q���݌j .&��fTq1��7���	���@\L0Ψ�b�yqF5̏3���K�gTq1��߸	8̏3����`~�Q����j .&�gTq1��8���	���@\L0?Ψ�bڱ���?O�{���m�ݏ�������4������1V�	Vj����Mx�&���JM��>ԄWӄ�X�	V}g��j���+5���\^]^[`�&X��o«o�k����MxMxm���`�w�	��	�-�R��.5�55�Vj�U��&��&���JM���G���M��-�A[�8m�mu5
���]�&�6�W��mͫ��M��-�A[�m�m�5AKm��<gn�DaM�R�5_ۆ�6�X��m�;��M4�-�A[��m�m�5AKm��:�6ܶ�ʚ��6hk=C��B���	Zj���e��M\�-�A[�K�p�(#�(%�&.3m�2�&.k��ڠ��>m�m�5AKm�ֺ�6ܶ�˚��6hk�Un��eM�R�����m�&h��Z׆�6qY��m��k�m���	Zj���{֦0�M\�-�A[�ok�m���	Zj���C׆�6qY��m�O�����+���l��̶�˚��6h���m�m�5AKm��}�p�&.k��ڠ��M��M\�-�A[��l�m���	Zj����ن�6qY��m�Ǵ	��M\�-�A[�cm�m���	Zj���+ۆ�6qY��m���m�&h�ں�on}I��S�6q�k��6qY��m�w��m�&h�ںtn��eM�R�u�6ܶ�˚��6h�~�m�m�5AKm��}ɛp���eM�R�u�6ܶ�˚��6h�>�m�m�5AKm�����p�&.k��ڠ�����M\�-�A[�h�m�]>m��&.�m�2�&.k��ڠ��A��M\�-�A[ϵh�m���	Zj����ц�6qY��m=g�	��M\�-�A[�Ki�m���	Zj����҆�6qY�t3Z��5����*��{��n���v�@^[`�y�U���Mxmѷn�{�v�@^o\��*��Xo�{�{�S^o\��Մ�Xo�{�v�@^[`�y�U�[Mx�q��{�W^[`�y��ۭym���W��5��Ƶ�jMxm���Wo�
�֛�^e�=�&0hq5A{�ޫ�3��p�(�jv���n���f�ܶ	����}��W�Er�&�j����W_a�m��	���^}�Y$�m°&ho�{�f�ܶ	Ś��}��W�Er�&k����W_a�m���	���^}�Y$�m²&ho�{�f���6qY����
�Hn��eM�޾��+�"�m�k�ݺ��+�"�m�5A{�ޫ�0��M\���{���,��6qY����
�Hn��eM�޾��+�"�m�5A{�ޫ�0��M\���{���,��6q�p���?N?߅d�4�Qu1�ʅ0�L>*;�<�)v]7�i��X1+b�A�x�� �!V�Jƨ$^�z	#_��0&��	#a�h�0"&��F��1*6��F��b�Q����`Tl1*��*vV�q��b�aR��N���sS������e��C����'����ĲrڛXVN;��i_bY9�J,+�=��:�x1�=����`�{>���(�|V�3������g���Y��cT|>�����|V�3�Q����g���Yo�Ũ4����F��b�Q�Ũ�bTl1*�;��F��b�cT�0*v;��F��b�Q�Ǩ�cT�1*����b�Q�Ǩ�cT�1*��F���Qq �O`T0*��#F���QqĨ8bT1*��e6��#F���Qq¨8aT�0*N'��F�	�Z�Qq¨8cT�1*�g��3F���Qqƨ8����(�AyJ|hP�C�R��Р�e?4(��Az���@zF%�P�<T*��C%�P�<T:��#PB�@=����#PR�@Y=����#Pb�@�=����#Pr�@�=����#P��@>����#P��@Y>����#P��@�>����#P��@�>����#P@?����#Pҏ@Y?����#P�@�?����#P�@�?����#P�@@� 	�$P�@Y@�	�$P"�@�@�	�$P2�@�@�	�$PB�@A�	�$PR�@YA�	�$Pb�@�A�	�$Pr�@�A�	�4����(?h@�A�������������)��Yu:e�����4c���e�����dg�h*O��TG6�Mt��F�+�X:��MVz��r�9է����z3���9��S,�.\ξ����(R(�v�՜���Yw#�s,,+�X�M�)Vܨ�1��]gT�s�S�B1w��e��g����k���^Ͳr���7S$��l���/�2���F��b^�!F?�X9��d5MfR����lW�(iՍ�z�]���e���[7�ث��̢{�\t�s>�Na���e��T��'�u����{y��s���}�Ο�e��XVN�hL1����/V�3�w������lg\>"���'bY�<ѩbJ~r��Z���Ͻ�rg�͑L����XV��T:�&�b�T�TyӞH%=P�'M��XVN�ء���sк�ʐ����\W,q�i��s,}q�s�٦O���]��ͥC�y�sG�/�y��s�v�����|q��ioTǮL˦�=�����)�2RL��|�j���U7��k�<�shsL���wd˸��;�������VE���a�vҌwır>��B��`��S�����<1Q,G��K�wĲr�����U�z��<�<�*���/nCg��e�|l�1?fe�х]=��=��)�T������`���,+�c ����e�t�ɲr�
²r�²r�²r���SH������`�{^J�3�Q�y!)�F��e�<3���̀|0F���<3�׏��`T|^=�3�Q�y�(o�Ũ�Q9:N��%��K����fWf���`��#VgY�`9_�X9_�X9_�X9�M��5�9*��Җ�W�(,Ne2]���O�"����c������#?�Z��)����Tx�fo�1DcF�Ͳr���)/,+���n�Cp%��U.���d�
֕`US�ѧYV�#~����*�/���0P7g��y.V�ҧ��7����{��\�ʹǌsvV;�u���R2E>nr��1��٩�c�K��8�=ŎC�����֩y����x�caYa��YO~Ҋ�
�]]��ſ�l��&c-�e��3��B��KA�OSP�\|]���l��1���)�4��j��B��qTy�F���L,��^XV���4TiCr�MRɗ�`�R?�i�ײ���2m��u�譲��ryӽ(�����.ɲrާM_�B.�SBߗ~9�Q���8�>�}�c��{�0�'E�+�Ne��Iϥ�ػn�uo#	��s,~[��_>����ޏ���{�޾���ӧ�?�������7���� U.);1o~����&ѽ�޽�%E���ν��|�s��{3KFde=�{˞;~��eZ�ղ*Ia���;�3�q$�W]��Q<��	Zw^�T���-�5I�ə�Wq��^��)��J=k�
���^���Y�0���{y��n�80�e�>�5O#����!CKɨ�/�����$}z-�����撧�eW����M"7�n��vƛ��$��^�n'd���^Y�ʬ3��D���́*o�pAyy�
ɠX�6��vmxѭ���nW���*I��Ν��j�W���J�Ds�����,����I�,}�z�
=�+��x���:ɝ�����JȒ*���W,���Y�"�HxG+{w獁���x��]��Qmˀy>4o��Yd)B��H���_o�i�11��YvbF/���1�d��vh���ޥw�l�ި�˲�J�vn�,6�I�B���2�?��������]����/c�(~�� ����Vl5K1軽��#�A�������(�U�$* �L%�P����D��I�^}��ь��IQ����;���"ɭ��ֻk���0�t�
�n����8m�9�  ,���9/�^aao���G��8I���)w��d��h�z��^	�O���Bv�������a���?M�]�q�*�� ��u����A��B�y�B!�<š�~�Q9q���[R���o�"��Uy�׮" KX� �[����J\9"tA��o^��Ƅ(����-�t_���<�l���emu�o^@pߢ�X� ��.�U�M^��8����,5��1�[�6C���Yΐ����w�M�判e�r�j�CDߤ(Z�]-G$-��#�VJ#�
�|��i9%���cZ~�*j9 t1�����TS}<�J�� �֐�����x ��� �eט�"��n
�]��T��Z����(ɖ#BWf�����[�cP���1����T��c�3�c@kȏ�/?G)�!�����߆��c���z����χ����R�E��^(_S_�7$/ɗ�u/M���U�� f���N���|k}�e���������d��g��B��8^p�V������~f!G ��B�@�������n�	�7�a�ɗ�>�Mp�����y��@�+��  t�����)�y���}�/P
�7�O�?��}��}��|�����|�������ޏo���|�J]_�C�r�j�N�j�&.��x.���ˑ!BPL�^N yaqo�Ϯ&�Z���&B���p���<T��
+P��@E9(�	�[)D!6��c/�(�&���L�D�i���З�;�8�6���O)�}9:�HBXb'�/G�����Zȅ%v��r�����m��٨R OK W+��/��Jq ��x[�}9V��m�z�!ÖI�Ŭ�^�ݖI��җ�q����`:,��/�Jq |��b�}9"X�����m��!�Br�rʱ�[��Wn�~����Z�?��(8 �Tn�� �S����O�6
�?��(8 �TnC�9�?��(8 �TnC�]2�8 ����܆��!�q ���S����O�6
�?��(8 �Tn�� �S�}��TnC��8 ����܆��%�q ���S�]�p�� �S�r�V��q���P�J��-�¥6��(�8 |�����Kz�p�� p�a��j�o-yjR�(�rz1��[w����n�8Q��� Ej�����2�[(n�k21��쏛Р��R&(��K�	���p�D�S#6q\��D!6qR����7���b'(\���x��ClCW�pq�m���.���.�c=,�� ����.�7=,�� �������O�C�8 �� �� j �Tn�L�Ōh/�����Ê.�{5�g��m�ۚ�<��ara��a=������~<�.1ot���0��[��yѧX�F/b��p���1�$݀��]�SKk�BvWp��(��NC��*���piW��L�=Qg�=>.��
ߝ�}��
��pq� tz�:��:E���piW��Lg ������v���O��G��Kk���O`:X�X|Ʒڧi����%~0��%���kz�!6` 4BB#\���Y�F�ؠ�6 b(E�5/��YM��`��X� 6XX�	s�=�+@G7k�R��a#B#$4wDs��j�	���L�bCB#$4�Es�g�	�����C0BB#�yv�9:�#$4�Z#��Ԁa�o@s��b�	���f�9��FHh���t�1��0�Z������YS�q
!��j#4��8����'����tز4����<�O������z�.DA�-`��FXwlBs�[�	���6������Q�O�/FX�L������b�	��nX��ŀa�l�!:�#$4ºQ�CtFHh�u�;4������}h�a!����:t�FHh�ucD4�����릎h�a!��)���-`��FX7�Ds����:Nq�8š�0BB#����9D�)`��FX7`Es��S�	��n����a���!:N#$4ºi/�C��S�	��n8����a�,�!:N#$4º�3�Ct�FHh�u�j4��8�����h�q
!�^��p���J�0m �2�[<:l#$4����1�����B�Q���t��Q!�����tFHh�u�~4�'��nr�L�����p�)��`��x� ��.���m�/�8(��$�n��݃�����a����m���$����M�j��d�pO� ��w�ˠy�v�,���]o����m�'���c�p�k��wö��ۃ���w�>��ck����U��}��G��d�Tp��9]����C��^���fe�{���)BO���<��G0���7�{�A����m_a�!:v#�e�W�p�X�o�8�1��0�[6|�A�����_a�!:x#�e��W�p��X�o�8�1��0�[6|�A�`��l�>\�!:N#�e�@���h�q
�-�uDs��S�o�8�} ��:�ޮ�������޲��+b8D�-`���#�
������[�|�A��(��i�LT4��(�l[A+J�ܲ� �xW4��f�i�J���^a�����O�E3|���������]H�OSUӬ\��䣲�ͳ�b�u���,�ۯ� �������[a����7�_j}c����7�_}c����7�_��|�~��*��$�I*B����2$�I*D�*�H�hľP�D#U��*�H�h�J4R%�O��ՀT�V�D{�Dg��aPi,m�&��I;7E�
X��?�����������V��N�j�X�� ��A��G,@��f<R�
x�*<��Hux4+��*�hV�3 ��R%�
x�J<��H�x4+��*�hV�ӤJ�
�xX�*�J�h�J�R%Z��T�V�D'U��*љ�:��{�	�[*^S`O�S'թ���Iu�:�R�zZ�U��U��-�=��%��*&I��~�+�ĞT�>�����^Z?���=/!,�=����q�"H=u�N!�Z�:I�IE��:H=u�z�(��Q*�(f�
3J��s�(^v�*1J��JLR%&��T�I��$Ub�*1I���+�R%&��T�Y��,Ub�*1K���J�R%f��x1^�/^����x-^���y-^���5y-^���Uy-^��bMRDbMʓD�,�<M$��E�L�<U$��8YD�l��E$��8aD��SF$��8iD���F$��8qD���SG$��8yD����G$��8�D�9�&�I#rbM��D$N�8SD�T�sE$N�kҋ5�Ś��#�&�y�bMz�&�X�A�Iq��lH��� ��kR��!q��ę�jH��!q�����kH��!q��lH��!q҆�Y�mH��!q�ę�nH��!q����oH����Q&')w��.8�$2(Vl�(ǐ�Tђ�yaPR�Cy]t�����HK�zH�!2z]h�����NK*��8d��##�������������)��Yu:e�����4cw���'�����#�B���M��ܑ��F��I��u�¸�nGE,s|u��!���4%�s�O]1��9�f��l���,s�v|i��/�BS����l�^�)�ݜu7��B��Y�6��x�h�<&k�97*g̨r�����P�}Q�j0���~V����j��Y폾��f���������ޖ�j�Xk=�p����ѷ�d5MfR���"v��I�nuУ���w�*�Y�6
�w�9�֍!�**~�H\%��E�v�y����Q��m��qc,sU�;Nv ��䂲N�ݛb8�C�n��������ԯ��m<�N�8���a͎�S�i,Fz�9��]�e��{�:��7��8Y���Ú'�2��;2f�[���>BbJ~r��Z�a�Ͻ�rg�͑L��{�\��sk��޼Z��dT���G,B�D*�:?i�������9�6����4F����UY�}�<l0�u���\���
�����Yۗc.c��/���#����<��#ݗxdݎ�b��@��ʜ��T���:�ioTǮ�,��=ƴ����*X����H7Mn�e&T��U7��k�<�s(�t��X�nx���Ԯ��>��_}��*�����>�Y�������U�N��}8�~(��D��w}=f�g�t#��vv�@����<Pu�}y�y�UtQ_���~ݎb���;R�}���Y�ht�^������l�t��4�ý�X��������`��j�����M�8��̬����˘�������:<9��(�Q}%πT�GՕ<R�V�l|�3���IuyTg��SRaUY�H�yTc�3 �Y�����3��z����<{k�z��j֋�N���Ou��y�zn�$��]ON���8�ޗ�r2v,aH��]�OwS��ѶK��`��G�,N���{N���{N���{N��q����8G�;[Z����mũL�K��i<���hb�i�?���~���S�+M�Z��0����c�����Y�������Y��tsB=Y~�V�l�꒵*XWHM�ŭU;�'��mx���	���B֞�f�[/d�%,s��bo���0P7g��y.�ҕ��7����9�[Q�ge��x{Yq��j���:�ɏ*%St�&��[+�vo��t;�"�}����ǡ�CW{�S��zO%�>�Ƭ���֓��";�BvWW�uqC&�a�)��j�7ʲ�m���D�S�s�[�U��$(�~.N2[�u6�R����;i���>)��XG��2�YיXf��~��ͫi��2*������/��Х~6�����+ip������T�U�*��:{?P6M��n��G��G�u�T�����Me��8�O���I��������s����9�h���uc�{{tV��������v�ǻ��w��7���g��7�����TGXW�j��Ak���֡�z5Z~X�l��$���![�nK&o�p-y�%��䀖�͒oY�$ˢ��,1.��˚���W�ӿ/0E��˿8�Œ�YV��e�ZΦX���L���/�[���p���/�Pb��,ӆe�_��e`]�,Z6򵅯-|m�k_[��"����E�-��Smj�P[��"�����E�-bmk��P[[��"���H�E�-Rm�j�T[��"-o��H�E�-rm�k�\[��"���ȵE^^��.�p�ܠ����:	Z�jh��������Z�
�e�:z|�Kۋ .
�Hࢁ�.*��`�-B s���v�-b�E�ȁ=�"ZA�$h�ً𖶋,h�- E�H�m�"Z�A�<�]T��]B�Dh�-"�E%�Ȅ��"Z�B�"���"Z�B�\h�-��E1�H���"
����]tC�phQ-ҡE;�����"Z�C��ٖ���h�-"�EE�Ȉ�"$Z�D��(]z��vQ-r�EO��E�")Z4E��hQ�K7���/�2��̢+��ցw�)���~_��y��UN!�UNm�UN�˾K���(_�&�Q`rՀS�q�4�;�q��k2��	��g��įp������d�UN~�#z-F��'mx�-�Z�_ꌢʈ��u�{9kG���,�l6�lC�ފ�_�3F�}Հ���q�UN$yՀ�]���]����VF4t�\�˳%����|�>���\�.��?���ˉ%%��x�I�Ⱦ�p����b�5��Y-a'l��;p�u�8q����I9m�	혽�|�Gk8Qg�u1?bX�I8�c=;�0�[��e>Eux�.ש���]b���q��^�F�%�׾E��q�+tt����8���a�ݠ��V�\H����E��ɋ$Q��,�Y+>���Ƨ���6�5Y!�Zi'��� c�8{C
��)~��x��C�dw攮���o`w��͟����~�Ok�q���}�o_dɞ�̽���)��+�Fc���82�̉��^����G�����kt{��;!:{�3��0?;��o����̯�^��m�~��3��|���0���(�3E�#�H��q��!��7N�7�0?ϒ| ��7�0?=���NDceT�������^G ��E�7�1�8�|f���𾦔�g����_�J>�Z����_Ŋ��gL��)̏=��M�Փ����X9����
S�i��gm��g��D�L>�����}��8�Yc�~��$rѥ�ţWP����� �?0�gVѮ��i)�������G�J_��0k4{�*Z�������p���,f�lm.f:/z<�>N�u�|�xN�����V�����F��v�gfk4�|��D�n$��^0��RF��t2r{������[�c~�#�^s�fw�����k�5��=�7D�om�h�""^4�w:7^��u~/,�e�E�']��^#�Ը-a�.Țo-4� |&��q�����y颠O2)��MwF�w�	�x�u�5�I�0�����_h�k����_>�}���C-{�/�y�����>W���+�x�֗��%��d/��%�xɯ/��Kn})<^
�K��R\_J����R~��W��Z�A_�X�AO|Кz"�֌��c����-Z�EO�Кz"�֬�+����h�5/����<�bּ�/:Y�b�x1k^�/f͋y�Ŭy1O��5/����<�bּ�'^̚�ċ]�b�x�k^�/v͋�ҁּ�'^��ċ]�b�x�k^�/v͋}�Ůy�O��5/����=��ּ�'^ܚ�ċ[�➞ݭ��}q-k��/n͋{�ŭyqO��5/����?��׼�'^���ċ_��x�k^�ӳ����/�x͙�ůy�O��5/����e��>|�{6��8��}x��s*Y�Z�w��=�4�%��K���]Y���O����T��]~�O5VK���!~���߻ϵ��O�_�����������%��X��N �k������:�������^}�柺?�?�U}]��u?}|_��M��O������b���s���T.~����O��ӗ�{���O��7�����}�i��?=LG ��������H
�A���������wƿM��P*dV|S�1v��VE_^ktzP�6�J�-}t��B��>-����?}�>C�o�߾�x_�t�o�����K���w�����op������m������5�go��}x����o�׿7���y�����+C忕��군{)�^1v���o��[��Vi�U�oE���B��5o����v�]�owy};��A;��n�<c�ޛ����qzx���-=�wo��ݛO�c�<��wo�����q��4s��Y�S��y��'*�!v6>�a���O�����
���?~��Kہ�7#�j4���J�Г�a�]�q��^���?kg�	.�\�Q'�T7�F�bH9d��K�����O��5����9E��4�ƓS�\]���l���9\���|�����������'����Y.�;3�N�Ts���:����q��8�tEů���������9>��si��JJ���cSuR�'�&����_}��4=Ggk{�I����ʨ���_�P�3�����s�����8N�]u��ﺋ���:H������}�O����~i�������W�����_�������?���������iC\��?�~�)`iʱ���ٹ�k˿����n(|���.d��a�k�L��R�쬶#�a�-����4��W�b���4N�\�X^ϳ���R�M�Y9�zS��Xޢ79�1ı��X`�叿{�O����>M����߾���~�������������r�����0=Lo��|���O��/���������b������?v�?n�y�~������_�� ���a>/�YP���~���=~SW�����B�v7���h�?�������_�7�ξ�E&�9�?��_+�v���[�z~�c��?~��G�����{g]{���s�:Z���iO-E��lU�C�
ej:ֲű�y��9�e���ik�ƴ�@��S�C�d����1��U��t�����>�(��.�Z����*�O:q_�"^-�}$jQf�E�LG�K%(�T��<�����`|�t��c,eުܓo��UͰv7y�����?�}]f�9�eJo��(*����c��*���������7��T�������3z�������ϋ���^���������X77�o�֑r6�tm�3����0=�T0?R��믾"�����c����}y����;�����M����?�Պͭ���?���������.s�O��^���+��m�e��_�;��Ha�zB�+:�!z���*�����Ϋ��:]��;��9[�0��O���P����k������w΅D��29���ȃ�8��٘\��s}ұt[cfeBH�4�eUyM�yAkߝ��=���?|ޘi\br�󚶧�e^����xu1=[I*>Дw@�~�`[��T��ષ��]�As~�|E1hS^�l�c(���/�6�X";_Ĵ�ɗ�vC�,_-�W*���K9u=���@;׫d�7:��e���|�� d��;l	r�^�wƖ�o��[j�]���HtƖw�5ٱ�Ж�nI���w��O/��0�ڭ�|�S9��b����a����P	�t����U�\���W?xqٽh�~&����F����:������������o~���/�	x	iR�0.�G����$*9]��e�3�"��|-�KG/�q
�{�I���g�MڼXM/*�����ez��e﷮��#���w�(��Ȇ���臵�C?�]f���su��=���*��o��������<޵�GI|���p�0��X�U!CW�g�Lj�T����3^?e�}��+��� +LS��J�����E!�Q��2�|q�I��!ȵg�H�@�]\��C�qfY�y>7���wk	߿Y��tigt�p���)c�K�wA�Cr��(Z�����Q����fo��&����1�s��޹����P &g��������|%co����'9}�Q�7R����$�H���3�����P]��R��(5_�S]Ko"V�n�<��5�����c��E�_ҟ���{,�x�R���3�?Y�5�k�/Ja�%�YGl�_J..���"��LQ�M��ez���"�n�u�«���g��������������X컺LꌫI�=��V��q(u�������^_����jJWWS��꯯��?�Տc�����p}�?�j4-U�1��5=�#������������JWWS��������������U����Ɨ?������r���u��}TC,r*�����tţ�`���ؼ[l�Y�䲚5�z|JTip��������?kgj}�d�x�Z'�]�qU�]����z�[ll{k���e��r�X� i"587OCG����U��3]�<�'�X���\gt*uT�R����=����X5�=\=��4�����4�abU��C�s������*����d|s�-T��1L��V�C���eM|�j(l��e�+�A��^un(��E�Cy��Lz|T��6��S���X�1YU�إ�h���^�z�s�+�d�/M?S���������;?́�=U��bu��:E��w!�@�2	��0_��)]�#9���&��P:�T���~*�Hw~&���:�e�ˈ�(�����L:f���7��O`���E�K���kI���z�ї)��/��S�6��RzWF2�2�����m�����������s�w���o�&|��_���~����>g��6î%�1�/����<�XH~*�k��|,2�u�)æ�s����KЬ�Ę�=.:�bu�+�8�ڹ��6m������7�ˌJ���ג�PfF�$�XW�s�ͺ�j'��-#J�c�U�Y����ظ�?~^����$��#&���>��_��S��~!��}|�Iuh��%��]	�u-��%
�Co�ˊ�7[!�Cl�k%��K���&k"�c���	��r<}Q������/���%iw	��˥��Y�k���t$�ǫ&��W�����u�h�I~��3�pV�Zc��+�叏_��?�����#V��3,Uu�@u?3O%�M��:���/k�ɮ��_s�:��,�/n��Ui�Zd�#wi���f������^fFi�w�(�ߛ��j��B��oP����~Y.��K�[�)_/�6Y-�&_�{E�����UG�[Ɖb�RH�����d�Կ��0=_�ܹ����\]l.Er�g��Z~5v��O�?�7ǟj�	��PW?u-���S?qw/���+p�a�S�ő��.����2%D���.{�2ֺ��s�ٲ^ݺ�~{J�6���}�?�n��l]|��i1��/��������,�����gңv�[e����1	������Ƶ�����珻���������n�p�q���A?m���~h����[������=�v|8ez��v�w�q��,W��(ۢ1r�=��^,���T{��ü�_���R�۹.�=�g���/y��Ku�PW�{���{RWa�a�B����2�Ώ]''�ӈ]~�����������y{qO�~{���M��eÔ={�b�ē�-{�!��<��%��5�|=��u�[?T���/�A-�"ѻ��K�C�]��/ĝ߅ŞwO�Y���m�7���T�u��n�y��{��;�m�`|���G%�g��;�_�es��_6�}9�h����^�\�e��.����8t����҆7�ȶ~��5�~w5�m�`s���� ����1l�w[C���F���mu֍�mu���m����m����my���m9έw�ᇷ���=�_|�=�>����K�� ��y��I����[�ݺ�`s�ܿ���n�j{,ݠrs(e�����P���g[C*��9�YI�%(��'v��pkʶ���9�&�~�1�۾9����[o��,?����`p��-�[ϲ��M7~Ⱦ�*ha1�/���k��z不�Q^�އ�l��`X���!6}F�Za�����!��i�8Sd�W"0��o�k����Ţ)����������jv̿�0(� ``���\������,b� �8�[@8�@0����q��À�B0�; 8�@8���օO�k�?�;||��'����;���� ̚W�`���8(��pP��
?!�B�`_@�Y@���B�b��q�����'�R�U �c��! �] N�q��!��_B��.,�1 ��
��`'�8�Ɛ��
��d�8�� �*x6��� �B� �x.�~����]�>�=��ҐwD����B����� ��  Ÿo�Nc�D�! �t@�=C�S��D� 
� �!�>I��9|��з����L'��L6����l
⠐ �A�ĞE ����4=�p��حVˣ�&��a;����e��[Ũ׮ɜ�w�KBY���Z�w�e�6��À�P>�����2q�b�څ���w�gp��2�ĩ2i38�n�M�8��|��[i�p�T?���0T������aBom�tzѬ� â�*�~	%6~k�P�0)��S��`ǯ�`�9�qK	{�h�H&��D_u�.�l��v�ࡍc�G⺎�;K'����d���)��"7a�rڈp�:N�3�w��/�30y�Bz���I����qO��GlӷJ{�=�1�b��T|݀���x����+'���1#7:PD������0{YL��N�ѿ��F#�����Fg�Ѩ��|��_�T��F1[w��.����f�G��FF<a���7mg2�t�l����q���rb��D���&2t����ٌ��~l��1܏��V�+i6����=i�!5���sj�&��E�-���8��+E�}LD�����4���''	����$��?�:򽉝�G;#��@�f��%�}��:"�I�Ъ�I7L�wM��[7�'�@#�]�7���p2�W�l�v44����bڌNO���u��4��8-L/����(���ub�ĸ*b����o�P��?�W�1�D�Ì��M�������?�t?>��?Ҙ[ƥ������}�~�4����_�=��׈��o�����0����������O���E���J�w#��BY�����g������apӇ��$h��Tq�i���f~?���x�b�Q�w���O?��_��v�}x����{z���?���w>��q~>�i�j~?�����E�]
xwV�	]���qJ�2�}�^�۟Oy�s\�t�����?=��4q�vjKю&�9MDS��649�R�K�Sn2<�lbo\���0M�$�����B�sX��DaiR �Z���f��s��8�a�-�_��y��{Ey[��vioItS���$�
�5��p��h/���Y�0,�l��[���L��S�F�B�"�!R$_!E���R-/=-�`�%�����g'6A����m�ژ���W^[�+�fҔ�� 4J���2Q�W�l�b� (�`��o��C0�@�B~$�:��.T��9!�0���`��Jq�F:�m��1(�B�µbHU3�y�}�z閪G���l�<E�ya�xj~�]S+�/�2>M�䱻�j0p�"3cQY��yk4D}�?�_�Q�߇�w���������Ɣ�W2�&�2h�GLT.`�����2Kw��I�30�_�>oHy���J>6&��Rdk"n!y�m�d/ }G�E����a�(EA�������D�O�b�6�~�R�Q�YZ��������i5���4�+é	�آ����jjKb\�W��Vw���`ԝ�(h�\���a��<mC%U*�Qws������/	u��G�ɥ�w�ֆV���量V�i"z�����/p�G��YRnrĖĐ[yQ�a�g�g՝���+���p�X;�а���vN��IM*�YK�~���E�����4�������,�Cc�p�d[N������O^iصl��!9���/�<g�R&(����D{"�����x<��(:7����5�����0`�ċ>�
�z�gP��z�k����z�x�u��6���7,�we_��:�B�ڄ�5��֎�J#I'�V��ٸ�mUVVPDm�G ��"�JT\�}e�nw�"��n����l�ND$��<�`���K��\k�r��@Ԇ�-�X������c���"�y&�]V������������9�"As���}
�+�_ϛ��%����.��	K�����f�:l'�D��?=7D�r��Qe���kE���ڲ^��yɖ�pl8��
�ᮨ����\�lgw9�)}�/-�j�u/��RI���!�) Y�2�s�'��n���6���F�s7zR\������;��{��-� n�Y��bn9T��+<���s���5Ǝ^e=��䤗Z��^�Nt\�����J��ڐh���DC�8����[�l���D�R��"/�6'��W��-���W�Ƽ�a�,��>	�B��% �9j�Fٶ$�����Օ�:�W�x��X�g�G\,J����q�,�l���a�܍-)$qA;JGW���dkE��5��Q�{nd:@c�������J"�@8���^fm̊Q`7:�����G�{���:���G�n{�1���?v��I�^o|"��bҙ�#���hl7����aH���t�}7~S����*3Bi�7E-)�AX�z�mb�+ÚY�5����X.b�H�D)�I3
Xp(�����x�x%]�Ɓ��ɫ����t�g���˺�-+Uh2[T*'kSc�>'��NwR�(1�p����d�e�}(�[�ZE(������W,����Ua|����v]�ca���.���Q|�Ѓ�J�]�G�a��Ae��	○�۩��&����`�IN^Y�yeҐn`sИ����|��b��(oL��z��Fk�ͥ�X��� ���P�t��K�=Ũ�D���g)bQ�U������e� �dmv���Ύ8'������(�ơd�)��)v���H�
gWPv`˰�`�I���ZXS�� ({��!Q�f��I׹����,��zK�y����je��NmP�J*���*��;�O�+PdI�W�0l��99��=�N�ZE�Ɓr���8P���F����OG�\�#6P��(#�0��VO�#X8"�'Nyo��㋉2v}�$�/�zċ�*ѯra�4��z!/d�g0�Cqҍ�%���u0hܴQ;Z/j˞��j�tD9�İL��P�a�~/���-��y�����x�'l�h5Ɏ�:"�ܓ�u��KTΆqgʖ�
D�4E�[��� �R2T#֜/��a�Bl��k�3kk�Lm�5^Ԇ��xBm���*��8jQj!a�kl�RX��E��F����H�i��r�v�Pv���48�M����(��f	�`��Z=Y�S��a��Y1<���gΰ%��]�)��}���e� �E�+J5�^H�pW�/kCA��(��2�*
xZ�g��n3��07�Rݨ����+�/&���y��Rk������7�����cs��Lڇ'R���~r����U�f���k���+Y#�3}�a46�"c��)oX}�g
�Z����ƣ6¯'V�-%ND�o���\:����6zo���d�Ϧ�&~)48�ƙ�IA%�^Nj��9���Ij�6Ո.���_[��Z������*��׉4�f�����������:7楾!fZ����f�ֆP��!�����a&b�W����M��f��̴���<h�͙�x��q`���g�,TВx�֌xU����/�MV�O����r���OQ�b��I���P,\�,X/�j���F��6Ҵ܋�TJ*���\D�x�<��dj*��U;L	�7gU� ��di,�"c�Br�!hu�D@�8����JL��/��W�9�����H���yȩ<"7�#��*������O��۹�L�lj9Ы hr%ޤ9���j��J(��Ř���0F�*b��0�0����ft�U����֬�����0��㼱�榓>{G��g�k�C帢�1�@�V)��, ��KY��8���y�n�j��'��7��g14cC��H<M�|� M�*�*��'g��l�g#��ɭW�D��Ѓm:��\�;�����6LJ i�I�"�b�iJ�j��\c^\.���lR$F3�yH��v��ڐD-������^�a;�J9s#:�4��xO�{*��A� �4��{�9S�l�V���41��+��ݖ�g�r5F�M�	Gh �(�sϴi�'�� (���|j �[��2���a1M�r�L�0G�ps�^���4�Z��n�$NaW�xU�5�j�'I����,qF�"7�f���1�h �O�νk�9����t�]�~sxI_"���Xf�d�~�*O�݆n'U	���L|���P:�N3�WO �v-a2��ڀ2������G�ڎ_��=s�C`��~�8ӳ�\���"�2�5�&$,�]/H��~�����피��mC���`,3�vIJ wLnp��i�K�-�j�����ϣ��_�&/c�(��-p Q��Ya�mh��Q�7�� w�yQ�%�7 J&糽����~I
�^+�RxU�DGd��ȫ��g��
��s�\T���U����H�u	R�|���������F�蜩ku�U���_D�/76�0��$�0����=��˽�a��Qe���ƀ����L�L���ͫ��ݻ�����{���7�w����4�н��{��ï{�~���%0���ÿ������������{�����PK   ���Xyɜ��  �  /   images/110f4c69-ce42-4daf-8800-65b9db14e3fe.png�y�3���tQ����F���E'Z!����� !8D/�[⢝Nѻ��{��|g޿��wgv��}vv�_vgg6�P_�����DKS�:��� ��bJ*�����K�����������I:_5sߗ�N��0(F@@����[���^PAO�s��=c����q���W�AO�]{����s�|ǋ5���5$��/�}�6�av�B��0��Ѷ���*��� �mik��Tr���ArlIڥ�z�!��lS�I_������i�|�J��?��!�����"L�L�f�>M�8�~SP��v"p�_��b��*�i��:�����X*������#�F&~x������NG�2Jr3��?�P�sH�{�>7��<X�̠��A8po���k	l�ʸ�x�cu�����[o�Y|��r��q~>௳ .��P�m�^��H������e�/�����$��4i�80�o���j��C��ޒ�<�M0Н7!���[v\T���D��As  ����؎>��8;E*F�Z'�"�o��x+�G���Ǫ���8�i*7ls���Ef�;��&�f�o.)j(kX��㉉�4��`=M�¬�x�W��Z�Qj�5��.'%lNVi�����ZᏱZ>�O�.��鶭LP4�0��F�}�P{�����m�9��#e�I�NRۯї&G���k���ֈ�h�54�
��ܳ�=ӄNzۆI�<��ΰ �8�Ż&���B�/h�;ykm�|���ks�_T4�-:���Zt]:�U�QL��X�d�M�P"{L��<�8t=�º#�QR����{B�hh�-��j�>�
�V=��d����~�?}���Ԉ��˽���[PUS��H���,WkD |��k]��!��8ex�y!}:f� �TP�#�x��(�l��e.��9�.�G����qy���{�0�8�����y�VN� �t<x;:[_��E׫���O/(�����C ��/�D%��{�&���R�����Ȏ����l�	��q��9�g��0}�)���$+���<�����?��tl�3j�2�I'����ȭ�7�5zW��=��!HG=o�_��b-R������1ߧ?W�c?�&����l���'u��ٕi����QMrˏ�}�)8!�T�����_����������ƅ �fO����1���dG��
Y�jƁf�?
��"���F���3G����G��e�>2g-%�4����!�c��)��rB�Ƕ� �v��G��%G�a��PD�F�/�	̈́Xbz������?���-(�� O�vA��a�{�nq�iGᅂ�_�"m�j�$^�p!ZVgL���T������Nv[|�}NY��(�mFz�׃u�Ѝצ� >��,���svSBy�:�K����e���vx_�JX���k�|-�[��NZ$>����gR!;g��<��6�
���ei_(l�����9�LV3�֜2Q{�(�~[�蕇�Ld�"�gttE\ݞ���mS��bt;�f�&�P�c@NjB��aa~�y�&�����Q�X�
p���S�L�n\�f�3�E���s���'�쬨t�؛r�O�u�f�֩��	��t��:�Ȼ�V�����-��!:�	�P3Fo���I� ��cd 3�Q>��k54Kl�xg���sI�o	%������lJT�'����:�6Yd�7��e��|t-i"a9u��Z�������#�����_Y��W������P>�ɥ�פ}P�;�_)Tu����O;��Kw

%��,�%��yܔ����nH�ʇ=���Ҫ��p���O��,��Sf�F5��T��NOF��NKv22bh�p!q�ؓ�����I�%R�O��Mw��h;���i����Seͯ;� Hզ���Z��N��W�:iֱ��wy%�7q��>du)��b;a��3�y�0۞*�h�������`��V�}�0~��g�E��&�>�vR�_��=PΆ��W�4hiŦ�W��<�̿*�0��e��Vt����aG���.]Rdİ�p��b�]d����&O��U����@*��r��o��G���}~9͂T�.?�0�y��[�v�xc�>�sc�o;sӉa��1������6"?��[m���%�/��1�Xs:o��%a���2��D�w�~�S.Q[���?�=
�KE����� �$P�"j�8��v<~{dR�����j��l<1�T3�d��%~#�`>ߒ���IҙK�q�l�TS<֯x�po���\���׀l�ʡ��D���
R��A|2�jB<�τRX���� 1Rc��R,�mq���@Y1����ݞ/o�?a��c�2�.Q�t{�D�-k.C[������U��.D�,Z�3��Ge����x�\i�OWZ�	|�#�b�@��^���%�,_t8�|]���t-%�1�y��V�qC����T��žډx?�}Y�[>;*nn?ˌW��̡TO����fOM_l3�eg�K,WddW[�~Q�EZ�����FS��,c���g���ɭ	#�F�c�k���-3�����S!n���T��11v�՚�
�T�����O�480��X���S�]�`�X�RU�6ŘF�&^u�	J��1_)�@��$Ĕc�t�P�^$�%ETZ2�O��E�`�iN?$�֖f\Ծ��n�������Xd�hO����!�=�֊B� �>;�2������&M��4�J�
�4n���d)ЧO[����7]�$��tO28��@<FӦ�,&u�������DӺ��F��*?��#��ٌ�%f}ƚ����G�垛�@��pi(���L����@ӀT����5+�mA�ؗ��"t�RCR�o�1�n�Օ���A��_��ӵ���}i.(��M��`ܖ�	�ʦ�S��N�Ԩ��X@��r�ݨ�+|��mg��&'|�D�����l�LW�h�_ז�+&�`�C��gx�;�H��ӥ�v�~�L���k�x0j��8"��>�����;s��,	�w�ѫ9L�vE;��c���n-M�g�O�#�@�k�r�_�φ��1���w�/�~��N���S�f�u���X��[��N��%�DjK�r��9����� C�R��xtMM�Jfm#^��1/\�n�
�Η�jra�\h�1u�F=��O��9
�ʄ��h���~�>os�߫~�'Fw��D�����}\&eE�Ϳ
B%�ڰgF�F�j4���J7����s��sY3/����]��@)_r�T�Ǧ"�7��+`�R���dǚ�$[Tt�II{�\���Æ��n�n��q�^.�E0G���#��u���"z$1�p�а=��-Tf
�v$�&*VKN��Ɛׯg̋��ʹ�o��b�Y���������:K$��@t���P��E��h�+��,� ��P��z"5R�dEm�^�|����;�Io�G�&T�%7k�rĩs��^���j|!p۫��!�`Dn�f�%D'Ѹ����v�	w�� ��o��r�� FT
���7TTj;�@+	9��c�<ϟl��V�W*��U�����M�F���|o���6�b#���T��htl쮏�����2�`@9���<D�U���+o)�b�r��2pV������D^�O%��.�W]�����V�XDu#la���|k�Mr�����j�sG������P@�g�'#[�D��sWR tO�y���d��
�M�Ϗ��(���$+7�i���DmNß#_ah�o�~��h�c`8%���s��?�X�*���	�6�_~SxX�9>ZD(V�J�
�z�`6d!hN_�0�z_"*�� ��#�僖e��
󜳨���Q���C�k�'k�A�N�m8i�����QAW���V�ҷPH �@�\�Z�����v��a<�,A��T�I	h��߸V�87� �:M��N��͹Ji<|�kމ������sI̺��lE�����h,?�ܗ�Ӓ�m�?��t��a�!w�rJŀ�8��Kt�B�A䇋��x/�j�	L%kb}��/# _�7�օi�*[Z�� ���6����辧���������w�맛ʭ ���K11 G�M��G�2���O�Av���Ozy�8�l�\�z�Z~c4`&Tl���/Hs�^*�5xw��R�т���[Ű�n�-6�e�!�Y����z�a��NͰ�A��&��a��-���ZOR�;0�$n1��-��L��!^�)s��b�4�������Ϥ���`)�9z��k���8��⭍���
M��(��_}�ȅ�/OG;$�]����*>R��s
���1�ثq��(߬�SϿ��|���Q���<�T��dǡN�v���O�xQ���n�Y	cx_��utd������ϑ����|�#nd»�����b����r�Fs����J,�WV�v�������fs������f��n�{z���jꂕ�.񾾘Q"j
Z��d*4Sm"J9�[����>�zӜ2�]�R�S_�|��n�I7M$�{�(�M#��X�����]�T�ک��1�UP/t��&��^P3)�%Σ�~��~Y�.e�I���a���|��h�׉s�,� �̅{T!fg���|<����vC�4^y-����@���#1�1z&L�-ZH�<�x�TŽ�����#^h�����Ogs�;Ӫ�Ѷ}��f �CXmos��7�Jk� ��3u��r_�/gz����@�j��s6/�1��^~s�bٷ߿n1x�ɚH�c���$"����N��r�=�.�mYQ@f�lt,=��z��pm�(�x^�*�q�sG��<�Xϑ^zv'|4�+�[��-5����e[HaZ�E���)�*H1�LXpND~A%}�"�H�.u���]�����([��aT䝌�y,4q�@F�m!���<e �S>�=��c��Ml���p�p��~���Ώ�٧ѽA_���"�:'6h"7��]��>�����)�Y,��!x��E���2D�C |�3�������}3bFꢌ
Y]�p�qJh7gC�ʳL�2J��>2$Qk�7��*����V�݉5��	G\N)����p�rU�/��.,g��t��yM���n������Ȇ�
�kp��T(�MRS����+��jo�z'����"?4]��%��Y��N� �a�����}3İ���p�Nd��]�AH�fԋ��p���T�T�������C��Y��F��e�9Õ-a97�����|���ß�p��#n)y �d"uO��R��g�q��اv�_*�_��J/y�k��+�Y
���H��P��'ݞw%������զ<~qhzqzǋXÒ�j�R/�A�W�۔3�x����Wb#K&W����ښ��#L݌�ԛ1d:0�Ov����l'ں���s���g�eM���{4�?�'��Gڅ|P�%��s���T�_�V+�g�-��4�*�q-�8�{��s~l����R�jv\��y���;럘g��|�XZ���z����Cqfo��+�eG5��ځR���K>�m�Ic����_��P<����~�w}����B77�2&5�{���2SY�ONp��Yp�4����VI8Yd�T��Cq��I��1I�� ���ӭ����m 4�(�J3;Ml��o^� YMz����*~[�1���Y���b<o�wZ%�<Î�o�u�󪴩71��tsmO��$ٲ�U�8����\x�b�cWl<��T"T�����+R��"�]&i<���-a�ŮՕ��U��3���`�`�P��8�\
j6�����o���4���S�.�SƌK0���~��/q�>w
�q��I�@�7�y0=~��X�����i5=�%MI�P^���=��Za=�~�����dk`�Q^��$����ft2#/T��_���ihD�<�����y
[,�������T��o��sm2�b�#_^�l�ݞ���U���=���|���3�&���B�H���ľ���':���j�M�����~����k=�Ĝ�Xkt��������̈́��������a��K��On7�6�ӡZ��:s��D�=���������m�A�R3�{�Ղd@d��"����O�!|JY��6����(}�F՝����C�Q~�2j��z.06��A�o@�$^,������t'��Qw�X�^zY#s�;{t7�y�'��s��H��VʗlHEXJ4�-�O���jO�?P�_!Z�%[T!<z��VQ��.Y79��$��{�٤Ԩ�Ι��K�*�*̖pf^�,= �g^�^�f��̜U"3Ъti���Km�B+�?��8�����3�j*$˧��C�ϰ�y�]�����*�'d�V���h�v�2�h�uY�p���H�B/��Y?-^�i��uf�B�q���*��ƽ��e��Λ�j?�]��nD#�K���d�=�W�L4���1��������td�����3���0m5��XB�$KU*���>^$�֫�2�æ���U���+�߻}k۞���w�~ó�O���Yq٨摆M��|������/b��i����8jL�X�)��0S�;4��6����f��|�D����V��7�Y�؟�kk���&m=��� ���� ��2�T��J��fQ�Blՠg'ٜe?��|gF��%���eo�2�W�$y�^���U��n婎J�d����N���|M��D)4P }���F���u����M�=���� s�LN�#F<�\h.��fY��>/��6����%J�+w����"G:Ӣi����,�Aj5����IO�$P`�o�DZE�:��q%�W����W����bV� ?��m���C�@�f��@����4�Jr�^iSt:�Y�X\+�)�]�s7���&W'�!c�I��^�|>��`oْ�J�S�?NQ-��I|��b�]5.��b�l�D��Y��U�w|�_�D+vE}�u70e&�C�3u�&O��ڙ�1f����5�`Z	�)}������
�u8��io�(P��1{m_	\p��*X�RTX���U��i���z�m7�t�:�5mSy qR�����,n�J��3{�X�Do[��p��6�|�j�P�Z@�8�CpVKL�9@��|i��F�jL+$D�^�݈�0����j�^+�?��1
?Q��<����,]���c���V[��/�!%f����Di��;���o����V/{@O�����e�����:؜	�����Z���?PK   ���X�䓶� � /   images/132fbcdf-34e4-44dc-827d-09a965026955.png�wT�Y�/��QgPA�H�%PP�tA@zE�&]���E��@�H��~����ݵ~޻�]�����9g����}�9񉸡�u�����赫 G�#'/:�f`�(���5�C�:t�1����z���k �w������)?3?COG?�m�u�p����� ���JS:�@�E\��/�{i SB����[�?���s�?���s�?���s�?�����
c����A��?���s�?���s�?���s�?���s�?1..l������c����DQ�;1����9[%����-���w}��.'��3;�\�/|���Wh��ж�w���t�i�%��_��������~�j��w����P��S��OZB�v�3r�r��E�8:`7�h֤���`b�\�o��{"?���s�?���s���Fq�� t�t�k��iWg%��ZQ���X���9�G���N�Z����谥#�鏀7z7�;��]n[�PQ蚭0B⏣��/���t��/wetiD\B2�Z�QF�:�+auY��f\�@�;j����+������'F��~ӣ�+�qͪɱ����E$��@k�]�R���.#}��J׽��L:�Ʌ�?/ZE(W�A�*�>��,�gT��.���V��`/�Y6�l���g��G4��乄��6K�E�k5�	/��u��]TfTz�MDڝ�==����D��T��y���
��=���]��|�	e�i�f���k�N�O2"����2hە�,^�S�Y@�&���2zf��K���y�ۻm�ʵ ���sm���Ȅ�WT�J�=~�	Jqi���.��g���r�u�&����&�+
2"��u�����}�۫����<g��:��sB��?����
�m݁k֢�97�����F����KؑQZ��v��6?QTj�M��	thf*k��}H���C��ߦ������^0����hKR��AKC{�{|]9��3j{4��������Ur�t[Uǣsml��o߿l<���"Vi<H���xb�lr>%G'�+�`]�h�O��6�rq�3
�gbxN�\��il� 8�Kb�iՎez�����N�]{�Ҕ�-I��m-�dTy<,5PF�ɹ�hX�o���md�^���s{ç��~��~�,|��; a�i�7#��ċ�SB��:�.b�vUrs��Um�c�ٹn��I4/"�Y���l��0��&�U�ptY�MY9����T����v{�ڞ�}O|�H']�qA?�.#)~�J�.}�n���F�H��H����S�u�O�}�)u��Ӫ8a��{��%����;����m��k��SK���ɺ�sYw0�������,DsUz�l%�
��ʒ��q�G�1釠��``��m}��Zz����k)%i�򣰺��;�M�u�*�/W����z���I%1ԭ`�@��y��䪧�7�SmƮ�u����u[���\��G�Ud�ב�ڞxݎ�4l��M屵����{�w�h,�b���Zzc؝]��	�#����Q:)��	��^d��Gv7�����I!�q
��>������ƞ� ��`0�Z�-��%���F��ڒd=�,Rm��WvG�A
M?W����O��/�;����-U� �����x����ǲ�^ 7%b)޷R{:r]<��N_ ^�}a���� ����Xw��>Մ׌��2I΁/]X1"g�2���@΀�jU�ۄK�"�l��Urn4�&(�&���/V�����K�[�����7��>��D���B븹C&�/�٦(ԢO1jk����P7��Z���봵IN�����v�:I������mEZ5�=�3�b2�߃��g��p�����Hp?M:��9����v��;b��Qw�Rz�D�,c�J����wF5�z�sʪFW�}�ޢ2z���`�̬�J4Z�(�2�r<.�&��K \R���>u����is��U���O��J� ���Jޱ������!<o�KVI��\�9���/�1UF{Z���=-1"�)�H���h�P�F(�ȥ�L	lB�i�d�bՑЂ)��1����#��~r�����5s�/L*�$�}YI��l̵Q߀I�o�4�2>��IXjھ���x����p4��᲼���$$��7���i���s��\h�o���ڤDBC�ս�d�u��u"Q��4(�_#�U�4���˺��2O�s�A��V���ᗛ݇#d��+l3���pC��̮sc2TE68�Iq�BD_@e�Y��I����-�@�H/��
s��7�~1]��s%��d23�)ol�v�֏��)"f�l�o��3��������jD��Q~C�i#��#�Z�4���������F0�G�1cط��6����VeX�;��>��>fy��Z�v���|¹���7�d����#�
��d=�2��~ߵ�Ξ��L�U��5���O�����ۇ+���#v-�TM�/L�&�V��ѥ�޷tB���[�mh�9��V���D����\��|D��v�X'~�1�πY ���)����� ]q?�Ӕ�����<�6)�xz������Z��UlQHG�y�j���� �G �IH�/�
��5�@��b"M/y����7M���a}<g�VY=7_7�`���&�b>`��e�P~�Cy�lm.]}��K]�}6Pt�V��"#筬vr�;�\���T�UȜ�� ��C;H���T���r઴fQ�js��&�V��y�e�-�G�`d�H�l��8
N-ib�����pK���S�Sݳ<y��mo�u�� �LN����2m�d��4�WR�w�<�azcc+���gz���u������V�e����.9xy��u��A-�&?U�U��j{(r�D^Nx���f�7�$���u�LȠ.�~㘱���ҽ<�Cg���'B�^Zz�;�=���S���E�U�A�O��*�Jn��<��a�?�ܐ? 㿯�V0��kq=:Sr95���h��-nԘ>^6����:�J���4G�����%�u<���
Y'�=޳F�u:�z���%���U)[�/�{�*���V|��>�4�e3Rrx�K������j1| TDH��dx�+XfP*3M�,X (�`+�2$ X�f+��pE�zf �������Z 6�xx)������A|�[JUN]�.?ʯ�3�>쏣ו<�p�v?;�c�dI��U�Cbg�L�����1�Q��3;��]�+�_�],`�;ژ�Ņ)pu"�E{P���j���5~4��GѿC�A=:r�q�t7dwz���{�E�ȸ����<��_-�Лo��׏%�4��8mD���>��{%�ш$Id�[�eYk0�m猧d;�t;B*��>[y�-��rD��[�ab:˟�ܨ��|�x#pu7������}��m��=�5�Y�
���|f��5<�YL�L��TbA������u���E�I�U�A�9��w�SlM�3wI�����L��������S��qU�ɞ��ۛ�x�L0O��T����}j#)ֽ�`�:N�ҵ(��\5��Y��um�=�"�I��J�|ro.{�"4�
rI}�����ux�Ln���[�q��g���/�u��\I��ғVY�Q���K�!w�2�yre\X��'���B�*d����"����ȼ�*!F�AΨ�8�B��鹻z�G�M;萉_���!��OL�������}��3���)0�Γ+gA<5����%�X=b��C��`��лk��=���[c��{��އ�X����f\O����~�Q�����0aru�*�f� N$�\.[zh�p�5��˫�E�Q��
�t�Ū�p�o���s�q�~��5N]{�Ŋx���b�ߢ�y��<��dԣ�j�_�G�������a�R�}�$c���5gD����������#;{�;���a�R\�o蕱��9����)�BBҏ$+���D�1�!�ĝ�8��T�1��|�Y+x3
��65���o@<\��,�0U�a�kJȔ��?�u���XTG�N��{m��
0ZH����U�6�Y�պ���&����b�&��\����y�y5����e"N2gK� k��0�xPҩ�/��]k�WYn�]��@m�E�^]ꍪ�~�Y�frF鄩�p��0&�;��{��ڸ����W8���6�R���bb�:�P�#6U��ms$A(N�o�6(nU���[{��&�<{�pV�3��W��$A�:' �0G�L��Ě� ����<��U;�6����z�d1N�8������A�ʃr�;1��s��E$|rMu�7W�y��P=������O�X��q�Kυ�'-��#�{�x�$��c���=M�b��MP�Flv����������ݬ����`]���'�Ω�s�V+D�5T�v���^��f����j%m����f�� �A�|>Ӿ��L���d��L��v" ���r��,_�f�Z��?O|��j���]z�����<�������w�!������n#�05��lo���6Q�^ǿ\xsP��^�I�4��xc�UG�A3�O�dݹj%�/���`�������(����ҕE��v�}��*��s�m��`���wz�/'^�N�!�p65G�˝��Fj_��s�E��w��ǫ���Q`�*e�r�>L@��VE�A�θS.��&��P �]���LT�e�Y8��O�)�I������8[}��,�Q6�.���.t��.&e}//�l��"��]5�	ZSIE"F�����D̨r�N̎/2��I%�"4��+]���c�Sv|�(0�ۏ5�U�M�ߦ�x��q��4��C�,��uEQ�x�&�¿�$V�&ۖ(�0Q��)U^��Fa��4�Tgu+���sC��ͳČ$5�Y`dY�|���U.{���X0�1�1�>�2�/zi��xl�I�M��G��Mh �_�\VG�,�D3ކx���ƣ�0����ZI?�'��J������F��Ѷ������իn��A]�E�4��j go�\�H:93yBBT�7��Zn��Pha#1�>���L�j(�*x��ڌ'��+TEQҹ��Uв����{-��0���g�m�O@̖,T���mE,=5�C6�(b ĉ�E��
��L��T�R?��M��V�|3��I��M\�UПZ�iTF�1��1�1^�'h�CZGl{e�,�1��,���^�d8 �u�A�$����N�G�αCl�ɮ��Sv?����˙�g�A�NX4�]���o�!��쌢�wYA������&��V~�܍�Q��`JϏ�nG���=#�lf�ٴ¶c�`w�X��� ��x�ӥ�<A�KOC��x�@,��#�s�vO��!�c�(V���r>����}� \U�;��d������j˾x�^:nv�xN���i�Gb�n�p&=2�}�(.�!7�����[ ���W%��!��zr��D��!��lm��Z�rr<Q�?��B����#���o��+�[�nA�}!�7@��b�>~�/mR��쵫������s�y���_�`-8à>��q�V����q���2����g�r�n>|��f����Ĺ!�BB�cm�	3r��kiǞ�\$��e���/�.*�1`TغJ}u|�Qa@�y?�̛��Y���� 2�F��|O�"�C��BRa�׾6X�aF9�oV��B������Ч��	��4��<T���W.��Z"D��\y�������ƍ߇�i��#Jz;�!4���h�}��E9��I"��
G}x����<�E��g,�0���A��
��.�SE������
�A�l�}�6g��ةS�uk��>�ghi�=+������>��k��c��|�Y��1#n��8��&�N�<<Oj�CC+9�+K�WXᜱ���R���>A}�B�<k^�W�qW�4$���'P��B�a7�q·[�A2<�����VSѐ��z�B[�V2{sȢ���|�n!���p��)/&���ΑU�W���w�6��_u�E��]�\���O	����)�-���I�B�y�́_sԮF��)5_���9��ܢV��sͼ2��˖�U��U�>��dX?9S�����F *���'��:
lg!;눻����G�B�������W���쾿���H�sV�A�/�o�Q���MI�=����J!�tWl�U������F��&�y�A�NB:��%�Tf�#��5�-"�����^��_��z���@����!l�F�'�(�X�K�1*��ދ��dN=z�p}�$wE��G�n��+��- ��0	�=��2j�Z,*�-z`�	ic�hzf��R�����om��^�����Q��=��8F��$bxE5+H�#*i��1���7o,��޴��s�6��]�ƻ�Wn铲���U;� �e@��-�͌u���(���ֱK��v�LV,rQ�rGE�$[	��<�7�k����N�ċ�myxn�.r��/b�6
rm��h�{I��'����|���W��%��}N)X��o��P�z��X-�:�1}���{�����A�iH�	��km�{���t�M�^A�D��A
��QNb�DO��Q<2������~I�����g�7��P_�N���E��x>���@i1��~:J�BU>��K�\.�(�"��ē|e�^c���@�� dS������4�3�{�'�<k��=/�>$Z�AQ�-������GĨ����P(������=�$���9V�qp�,�y���o~�]�)=����	 �ziC���u�7����J�~�JUE\M�T��Dq*j�^ �~�N��T�5�L���O��1+K|[�x�s:�Dm�My;�W�����~;��	�zO�Ჺ����!�2�bc(Fq]�<b���v��*!#_�ַ�҈%��]P> �E3h�MT�
^8��ӳ�~�6g'�#\��\g#�7������v1��������\�<SG�_[ۏvx��J���d7���_� 4lご4��.$��l��Wn���OhŜ��[V���a��gM
t2���%S�ĬF�A� ��Bo�|�[�{GN��߾i�~��2�I��_�"Q�N��}���^&uf@�W����� d�"�i�,���z��ؙ9N톀,�`�mF������I����o��l�4Tx��W1�M���?Cn��W�7����;z���T�glŜtH�ߝ��'C�!��?TP��C���������"
)<۶�1���4����y�^�v�yw~�t�ze�f�5�{!�Aslgc-�Ge���@)�ϡ-��z��*��8R�����Q9��[�Q������L�K��W�%u��}18��v@ա�hg��}{{�GyF�Q�Ql���7pc>��Z?Z���������(�\�|��$���5������wh�G6pg1P��8�c�?'�u[=�J9{��L	��I�-���ݭ��?rk{��܃nھ�X����@P�p#���޳SB�&�ˤU8�ؒ�?`=���Z�$�8F�|�=�⋠���	-Y����у�^���}$�u�ۊyj��yx-�`�Q���Lp�Q\*��@��aЄ��t?���jp��DNj$�LqV3,9�R���O݆��;3q�(��5������n�x�b:�!$�a���26����(J總,�=
�0'�ϋ���!+�TRPPWJ/�>��T�L��m�~@���jnI�݅{�4&D��
��ܔ��4�������$À�"}��q(� TAG��4��K˪���p���A,�o�\j���|�D/?�3���y��@>`��L�9�K+��W��Դ虬87�ڑI3�a����$}��
E�,�
o۷xŊ}�@F�X$@E.\��rf���R*�1���x���>���\�L�����RSM�Q���yOX����C]DlvL�M�s;���cW�p(�ݞ>,Bw�^�?=��+��%d��}ˠW�Z��k��Qx�3� ��o$U\]���u��l'/�D����VP*q�`�k�Z�ݓ��V���i�D��C�N,GJ����)����4��Z�ɏ.\�2H�j��I�.�S��h��5��M����ʃ�A�)s���읔��_��q�uC��q�8w���.xm[)pm�bpm�I]�~=w0jZ�t��e���`���A��A��~T�>��j
$�mYМ4#p�?�#rg��'��Yh�;Hj�eWd��w���W
6�{Rs�[�`?�AMy�#:6�lyB��� q�ի��}_��6�=܉���j+)��� �L坏����j�)ۼ���3;��Y��I��7$o��������ZicD �l���ksv���VjP��l��&F���pd�&AM��m���-MG��*�̏��B��N�v��F�9�M�C�	�#�~2�����CsH��Q>3b�PڎSna*LY���;ڮۂ���H���"��O���#���/��K�Y���*��P�W>���k��m}iCkH0\r���	w�:��ua�3`��k�w1�`�~�M�U���ـ�}�!��;�`9����Pw^�X7�[�LU׶���v�cKѽ�a����!tf�NYL#Yv�	Du��#�y����̭�_mF�`���
����ka�ƥ�W��	��dj���T���ؤ\�[��\�W��]Q��תv���ci�wh�!�@Y�d�B��LU���5Ņq��Pw�Z�ж��^���a.�*%� �Z���rߑ�n�����_l�?��x�x������o��b��u4{Z���v�����αQ�T����WN��W�&���ɛ��I^۷Ѽ�Z������OT@]$��[��0��K5�@a���ۂ[ƀ�v�0K�F�Ԙ��Ǜ���˗�H��Ru��s��DH��/�DR���9�F��jS�A�&Md�f{U��f�M�B@;B���؄܌<5�/���:�+Bѳ�B͙�zaB(&Bf�F�#gԅO4��Ze�]{�n�eM9N�ʁ=U=�uKc@,#>�n�l�H:����f�Ǩq	4m��>�g���=��K�yG�^�~eM���1��Y�w����^��7x��V�&�����'#�8��=������rSQTQ�6hs�eʓ�\m�����gi�=֜~Ec_c+^!C�݄��?S1�""1����U��l"� ��/ w��6��Kk��1\.�����%� ��#�j�#72�C|'��l�����M�-w"������7�0�����h�#���>_cc�7+�����T<��0կp���l��^�6ȼ�:�r��|�m��x)����{U�;ӗÌ�Ƃ��vJ$��ڟFo"�¹�n��H�[��`��S�@;��$M���Y�V3�cY^�|�X2�w��wْ��;�p;F��jo}M,2x��FuǺ�w�@�=<��Su|j2��R�M_A����Y����$e�%�/9v�6\<9���8��@�m�tY��2̺� xmGvGi�L�J$W�[�����6���&���Q��Anv}�S�pb�8m{`rO��\:�N$�nT?����w�i	�n7�O1��"�;h;�΅~5�>jj�[įJ�(��J��e�/��}ȓ��=nAC����).�wd�V���,�\ś�������4D�p�vB��аo?̟k ~1M�&
65c��C\@��K�.�R�郹�,1�H�r`F��J�,�O�����G���U3wgiB�L�v�D��\"P/�6��%�f7Sm��+Ӝ)��|�g&��qKި"L�?��4���u��r�>T�lu�b�У��=���WoS���M_�F/��KH���җ�6$���(`��a%#$�Sc��[;t���9�~E\1q�b��'�0����@�e��|c#�i�+�]k}����j��s�h�W��&�@�v9|��J�֜��P�gZ���V1[�٬#'}�G���R��}��ؘ~5�mȚcJC�<����9������b�~~-*������2�5���K�*c�X�=Z�R��س���3�����^�Q��"J�o��sV�V�b�����dB�e��_��ձ��,P�ٝ�T����w�����kaJbm�ѱA]i���hK��ظI~y��G��&0$�!ɤ�X���9��d|@�Mu�3��0��%�@�Ѐ���X��a�	�&����N�we��M8k��~�<
�PYj;������?��t�ϱ(!�}�H�4 l��{�x���Y`�j�;�=��C�<��wd���&�{�n���POM%6�#��q�>�0#1#4���:��!�X�0U|+�Lo���A��3���Σ"��3=�t�z� _ꔭ�\�;���L��k�3{��d%��,����@p�U��}k����w� ��o.!��8��ɦw`Zh��wؗ���W:���}�^����z�?���@��MŁ�I^2���P<^�IcB9��������w�"_�S!'S�8�7�����P��
�EO��\��xbuݰ+��qߚ��;�<聲[�w�VS���{��� �N�f�@Ƨ��Eu��qb��T-ǴD�݁�$1����T3c��!�V_�:t���4�c؟�9`��ÖlObN=/�5g�>�U�6�Č�Ȼ[R�^f�� �.���0�{�=�(A��Q��k}{XkN1��X��`��NU��h��0Y�f���]=��y��5GoM������x�
.�t��F�v��.�F���� �e)z@��\�&��ʼ�}'7-qv�)������*�u(;չ*7gh�AM.E�!-��Q}Zި���e޳;�Y,�۴ẽ�֋����|�}{N"J�7��-u��T��iO����q�u�96c��{�|��
�N�AHk��m�^�T�X�'���x�����0�"�M�a=���Wvk����'�q�k����Q�:�C��.���nh��zu~��z�z��h: �-[C��6��N�ǻ��a�`�l�_Ā�q�:���2�i�F�Y�K:�Z��S�4�6�_E����&W�k]��z��I���g��׭��[�`�=T
l;�g���֓5���ꤍ��r����n���4vٛʦ&��*4c���q[:K��/�G滑8�7�M��=���'�m7�K�A&o�Lu�I�S�o�4���&���(�J�r6���W��o�?v��@��iWY���$�Wty^���eo�/U ���@����Q�ٞpG�{�/&&���=[4G��\p*�p��1l�A�A_��2y�3�/շ����r�޳���������l��.�\�V@/��	����?�/���_�R�#�����'s��]�x��[? M�[U,�'�3�u3��&c�ga׹�j� ?�+y;G��_oR xg+����՞	���Cg.*�󒇛�,�i�1Vr!P��Js�>��^]ҫ�؟�ZC�[:�z]>�R�,�<t?�K�`��Q�^r�]��]N�N\���&%v8&���I:5��aw��Ƽ����fڑ��N�q����=��zN�|C��g��c��?ί���@��s8��~_x�n����kJFy��Z�3^��6@��S��U@��_l�%���.�l�m�-�=�l�	8#9g�lX�۱9���D�9S*�:LDx��2&��c\
 ы���35b-��`�iA��l��F�Y�:��}P�ܧw�G���ge����y���0\��7\EG��e�*�CP�罟��N�<��z�k�uOLӝg�a�P	�+��;�r�xE{�}�F>�xQ����$C��%?��l�g�Li��X���)w♴`�ܩT��/F�)�@�<�����ש y��w����ea�a~����
(����Nb*���v)\�~E/	H�ŭz��?�Ԡ���^��}���������^D&7_���>z�-�� ol��8Oy����}-�[�djGY�� �9�M�'�-�~_��Ě^�U�z�}�o����9I�ᾈ&T=
���/7��*��"n�!]-Y���/$v��
ޯ����i�f�ݐr�^��!t��<��T���2�j^oQ_����u��߮]}'$�w}���j�\�@+n�7��$�VM��'2�!~@6R1��Ȍ�r��b=���f��J��ә#�$�K�-4ݒ(ޗ�}l��؇4�o@Y����߷ �����A �Q2�>��#e�[G~O���<R��!��n��*�케�$p���W_�2��zƌb躪Dj�1������]Z��G�J�eX8͕��U�Ž���M�a�ཡ� �p"�i�^Rm<!�T�S^^%g>qs6(�U�K�8�ӡ
A�~���^�p���o�I+�A�
D����8?EDM�d�"Ԗ&�V�Ӯ�I��a}����-L �M�������f$qx����):��"Fف��j����o�7���K����#EOJz�sC1����q�P]|�$�l-�bB�����#�gX�%d{X���m,��~cw#(^)謱�nMl>�@���yT�S�H"\�ˏz�S�VÇ��KaX�*�t��`䮘_B���>�X�Ȕ�ں�~0��t>.�
mj�6͎+��B� 6��n���bf	�Wkj��L��pZ���&�[�u���*���p�m3m:�-���q�D.�d6�;]W}'}�ϥ�Q�)E�۬X�j�>^�G��G˘�p�@�+�ڬ���(����ΰ8:O�J���ĖL�y�JC��N�!�T��xQ���u���[l�A��O�C�%j�<�=����B(�R��l7�
���`�uf���\ bH8L��������I�r-Mȉ�*RPw���]��:��~\\t���/�^��zD��ފ�e��0��-*����۟>����9z/^��!~N��i�E6�����'�S�U��=�z���{|�p%����U�OMvU@	[���!�$���Q��]�[�{��biU������+�`�)���k�v�7��u_ؽk>Q��~�%_*yl|��a�ca����TG�577}�����-h��k�+���Q�jq?VY5ഝ����3`+�d*,y���,�[y��nN<��J]D��)�U_���� �~`�NU&�s՚�F@�z���������qS�� o�e��yJ[�*Jo��5fgO=��H*"CwR���� =^L�c����	6�Lxu� ��|��R1�b��'B<k���M��&����)����	�	"PO��~ rPγ�nO%h���VI�okq@E�g�ԟ��U`��*���L�xp��
�"i���HiA�a�Z"�ئ�ę���O�cZ��cgp��h��Ls��LT�R�2��vnI_���ǈ�܏{�� O�ߨ���\����o�ꘝ>���.��8��Rw8sJ��kj.u�5�*/��\_a˂_�=�?o��$�YC���w��lC�B��R{8�[�\�K���E�*�w���7 /��U3ơ&����0x]3�e�,C*۵ek�B��X&Ǻ/2��c���![Ҙ�3@-+zاK�-�_�#�~��
�/�i��73������gp\ԙ#��:��yb����(,�
j�L���y����%�@	��@��ˎ���2��}��.���?�j�j�˸
�8.�ߙ�ژT�/�ߘ�<P�������ŻN��	�-A�t�}�<��i>��tP�L���Y�ʾ~�2.�7�{��
�E0�V=��=Ӫ���/#�b�t�K3�1���N��?`@����z�D���$Ѱc���� ������c=�Ы����׏<������<��Z���c�;�2��!���� �u�Z#�ef5/W�`�m�'M�;�#bU���2��p��ѥD#�`/w�����~�ꈘ�>K=O�ݷ&m<�j���u��n~�����\�zt mp|���`"����1}�D�+2�/�Z��l_X=%^l�Lv]�&�}Ï*\aFj��ǎx&m��0�@�Y�Ws������&A�>�1�Ui/qs��Wb��UQ�s9-����}��Qf@�:��B����lA���2��͌�y��m�5;�z�޷�.��������ahm�y?#W������!�3�����T	�q�ά����i�Lu�|�h�3�c���U���M�?O��̔	{
}C�zu�s��ۂ����Mm!}(
�������uD?����\�����s�˙��{�,���:�XШ�}g��@APVN0�����մ�E�����<��R��GV

R�V~l�ϱ?�^���O)����l�<��:�����uKĵ�'��`�$��dr)�.��FID]�zP���LНC��/�\���"(gv�ٮ�f�o�S��A�:]V��;TrkZ�~��A�@mq�@���i������m�Ⱦ��yfMN�{S�U�Zd����V�%��`^���Z�Ic'w�����<,��^L���9Lb��쎑����(&�U@��e�io�!]n�ȱ6�(Gw��X�!b�)ڦ�xTTۨB����K��l\�/Z�o�q�nW� �l������&�,>����2��U�(�M)���?��{��xY>Gt?�̠%x*<����,�(J�R��+��oL���+Ø��c��wo�|,p(3Y��y3S¹d캣�=+��1����D�_��+�W��� 	����8��$bhF�v���aoj�_���y�I��ҕQ�X?f����;� ��R׶��������'�4�	o��6Kܻ�q�\���_��	a�k��6
��a�ʳ
��v��!��k7XD�2�y��P�İ.}4H�\�&��ˏQ�(֔89U�~-sM����M�`�x���Eu�L c{l��Qg�)�v��?!<'�)���*R�q�� �dwIp~�Pn���X�%�8�e�-�4�4�����&-��h�1�]�� ��t�3�ke�=�.���ϗ�k����m���@M��H�m/1��T!���>��Ie����3����u.Ļ�n-f3�J�:�ʼ7��0���1�8��g��.�h���Ȃ1(��J�ŧ�c��PA�Qǲe'���IƶZ���j�52� A�������xO��L�[� TPM�6����.�Q�e�}��v<�S��
^?vN���������8H$�L+}kbJ�Bf7cX�B�\l�J�3�����ȷ��M�ۯ��T�~P��T�1Y� �zo:V�8���v�~p Cf�;�>Р׏���$���p���jJ�5����I/P�{v,���^??Z�*u� �2բ�j��.�"3F��<s��F�<%���<z
k�8@gnX���XF�X�*�!sZ�퉙0WO�@��_�-�[2O�[�^��=r�+�m5݉y�>�<[�NGm��Z���VOn�+�$�G҅ 4R�VD|Ջ��o��ʄ�H�!�}���x2
$�O]���b�t%��׻�����!S���yB;8��OGϘ�p�Z�97t�h�ŵ>���!�2,����_�i�B.��틳/=Z�(d?�H6f�&�9Z��vo[�hL;2j0���Sb�vS�N�FG��X&��v�C������ e�R���'`�BE�;L��x�7�	r���~A�������F���MJz�Ci���(�'�,�=y��SW�0l����ۓ�RLY|u	�8�Yh���nf[�X�ڦ��
1�
��sUd:����E	��<���<Q1E'eM����h���}O�;)X@\1p�4j���AQ(� �YG��91�z�����Ў�H��7됆�H�:4x�> �ɱ�ڄ<C�տ EP�)� K�s󔸩VZ�[�)�#r���T�pӟw͝�P��Q*�W�
�#��o�����b��]jo!�̬��
��w�)k�G*r$�2��J��ǏQ�`s��!�?����������r�A����;�UA���<ٞq�A�x#��V�n��r�<�͖�mWF�
�L3n&j����
��
���R%���:Ef��J��ÿ�5�O�ɂ�]�q�@qZ^�:FIFW?��u��ILvC��M�߽V��;�#<W����I�N�"�z���})L�d�∃���s`��9�E�X]�C ����ՄDk�T����z���~<����J��Ob
-z�9�K���>S�ٟW!����a�6�<p���P�Ds6.)@Ԧ�٪�p4r�3 /�u�$��ؽGf�t�>�ws)�x�L�fy�A����wF�oѸm���N�F��ɇr�AL̎e�(oW���$��hpB���p��<�H{�ѿ4`�}����.x�?���-�Kѫ�/�m��v݁�?�5�4��Xގ��&L)5zW�`ypD��5*���L��su����BP��R�<x"L �x'��t��t�ٟ��(c:^��l�3[�}��;��uz+���4�$4��d�<�"�j��m�Y*g�{�9���<�(�����!��+�>��|%��8�Lz�j�P~�����&�:����ڋ��ֈh��̑�@1�C��.�I+����,�M"̰qS� }�Rt��U�����/��X}�̭��]�Y����xө3s���R�s��_ؙ=_s{��ʎ{{�����k�ɷ�)5aW�VQn�@ӥK���/M�X^c�Ŏno�j% �����6h&�=�j��j?�V��*�+/��n]r&O'oT�>δ)��5}Գ��2�NW����o�[q������.ϩ����')����M�e�Dt���_W�<�	���?8u��(0��T�I(���ԙ
�!:u�[M1�ߐ-��L�8J�׌rX����O��ob���P8�W�c��B��Y�>�	���7��@Z�������ax����� 7��\�Ce@%I�+�?p E���H�ItcV��U�/-MD4齾3�G[B�t{^ ,4&��A]�:n����y1\��ÌߗT�2K a#��;��hĘ�H��xU3�NR]̀�]�2�_��6m����M7�忸	��n֔��K�^�UC���@bZ}���9끨��J %�qE� ��gpYm�[A�zq�7�v� lۏ��~{�GE�7-���F|���]�������:�X��	+B��uI�e������뛽Y�.�R;�g�|�<Eu������ e0���NdJ���K�,[t�~��Ij�O��*��;�ܷ���g��F~`��8���6G��3:%�?9�l�g?%����{���'���#��ב�SL�M�__��xkd�YFh�]�9n��}i*L:�Nղ����t;���VJ��\�`ݻ�`�D^G�$k}�5?=c�cn�2$w7n��?r�c쯍��JQ鯩��E���Q/�!��%�1rtS��I����\��EL�K��r���\Q1(q�cH]T�פM�c ��|�nU_�*���Q�1Ǟwԧ]V��.sS.㴳�＆�ɞ�p8+��dE�+ O�ʶu����=a�:�i���4�����^3�5����\݃��w��Źz�����m����h�D3K�D����fy7�?EY1�]Ev�9Z����h]&Bp�H�/�QK�HE{��^�\Q3I(����`��f�C�N��ޝ;Zɲ��Dc޶ڼ��Y*|D��@b�4a�l8uى�6��������T�Σ�����ڠfV�f���@�zMm�z�<hs]��o����b�\d?޸?�C�Ό�.�qJ����ͭ�H& \�]�q�T���?�����&�L�s;t�l�?�����m��
�[���۷6cc�=���fhv4��������z�x���|���)KR�$%�%YO�%	!�d�'Df�t(E���c���5�0ʞe�����n0����>�������C3���}]������z�/
I�2@�◭(ݎ�פQ�۽���*�ȿ���f|-��[�V��Wo�R�3I,�I\��J�8�|�5�Wa�Y+�J��]���[�T� &:YRH���`7��n��H[������h<�n1�u��!��&z�}�����,f�?��V�u��C4���)k���J��d�������.����^{��gǪ��6�=����s��G�Ro�H[�ͪ
p�r^��P���r ' ��[/�#��.ژ�s�uc�B���Ǔl�A�up�:�Ԍ� _�m�q�XU�C�Ҏ�(�}���ϩ�����fV�P�I��a�!BUՙ���@���
!��\ۓ�c�o�ܙ��.9m�=��^�D���c�j����� ��&u�w."�W=���&��d�\�f]����G��Y��0.������F?*��Sk��]�wECx�;>>�Ґ�;"1!ٛ����9�+�VD�k�XgZjA�/t���d$����z����j����O�4@�A\�����8�5�Ur����@�@
2l:�*��(D_���:
�I����������j@ ����Q0���X]��I�E%�ox���3�p��8�۠m@<o�bPq͓Rv��Ǉ�[�#�"HlH M<l<������=r]C�rt�����a�L!ߟk{NU�pΌ6<qq1կ�M��I�N��ay����΀RQʧLX��;����2���\��-w)�?��'U�K�?0Rs���C�~�0P��$Di�+��L�Ҿ�TlU�� ���󠫘�P�	�drI�4E�[_��X ���B�qV��w�h�91�^o��l�fS9���S������*��<@+�7����s����ty�̥�� c��Q������ٲ��^ԥ���"N�0�<��xrU��t�}�����7+9��S���C���:�C�EM�v$�(�ٖe*\�)0��Â�hYYY�c������ID�pY�@��*%�m���jӱ�z���u�!.��k�̏w�y7�u���J:C���#��������z����&���a��i��������wUJ�=��mӍJI�gfc+���h���D���$�ښ���c����0�vPo9/{��[�y?cx��!�������L��b�J����vC��������/�������1K�s�į`�qBE��d���i��s&{[4?'ޅ��!Ấ�ib�@�n�.�r�Z�c�Nr0���~�����m��UNPC-m���-�(��L>�M4Ց�G��,Fuj3���<K���͸C��}"�lc�zI�`���T/����Q������L��⥖�۽�$+9G��0��ǾZ�h16�D.=�jϔ�t��K��Ѯ����L6�3Wl��t#��{V�3��!-D9�������(̄�PAa)�����˯ɥ'W;{�dw�.h
|���ht��-oxK��������50PB0��r��>-�?/7b�]�	�h�Ȣ�c�Hv�G�O�ٗ�6���T���q�O�q~f@%=�fLdA��G�	�7K�U,9��̍�׽ �S����6�z���d����6˝�="gc����yLZ���[�}>��#�/V
n�]_i�����h�p���^ �[�%ĉ�/JsH����	JVɰ�s%�{~
��L���=H3�Eή�a2���X]�҈�O��:�z��M�8�X�����y�6dOv�}�h�K]a���� ����M�/�FR���Q�'pu��J��J��uDD��U$-/ծ�7��1s���;�B g��B������!���_���{6��P�v5^ۉ�Px�K,K�8���ؕ�����.�yn'��T��H���_�C���Z����*X�WH(s{�^�֛�֩���̊R��24��<����}�����E�c���;]2������j���p5yX��y��|G���j�0�(W��e)�SF� �tKj���h��7 ��*m�%�C$L?Eo����\RX��g� 6]05卝���5�߷΃�<=��󥫫��(��RW�;��J��B?4��1���K��L��I��!��cL��ǌv�7:d��ʨڛIo���^"�=��)!��{�5@O�p%ۚ����]��T�XI݋ʀ��/WG��IV�+t���[�: �<��F��5ݩ�v�?x�ִ���[cϔL�N1>�E�����x��|� ����S��ҷ�S(��eHQԪ]n��?g�����_$��ٗ�J���|�z�#W,#7��i�O����7&sY�)���ߴ��2o��kl�
�^��b��mպq�Q�S��]�:���/їL�&��
��vO��6ٺ��"���'퓸�����Ih�I����}������{��`���3��w��Xt�pＡ����J�8Y��浦��{/OJj��Z��鈌P��4�.��/������9�Ō	O��2�VP��5r�0�j��|��Gk�9���7g��9E���aD*����1�d��Ȱ<���H����Zީ���m@Eu��+�'S�vڣ�j� �/�ڔ�\Is��@)�t�A��+1������be��=s������+�j�m	H�]<�ut�.�������χr���+̭�Z��H���q{6�8�漣��n���)���V����с�i� Z���z�<ڽ��
�`lѩ��s_�=x�}��*" ��F�OhiZ!u�G�j������\?�\~?�(�$reЖ��)W�'Ⱥg���$�����4و�W6��;j���l�i�N�`M�N��+ks��93�ӹ��I��F�m�s��SF�'T�)�pk�f�$� �R�p�dc�<�t�*D�*#"��i��㼑�E4�N�`o;��	 $Zi��H�0�[z���q����ߚ������9�%1GҸ�밬TI�ҰR9��)쨧,�S��f���f�91>z�yiB��7���9O�w����]u"�/>i�c�G�Ba6Z��d�������.�������e���L��Wh6;G�U`us��g+c��YG��k���ƑS��,TOH;�%�)���e�F$�A�P7�oM�Rk*-���k�����
;��XDA{Z��Zx���3;���EJy�	T�����С��E�*���3��IV��ӡ{��>|�λر���h٭�:�z��Ӫܾ��V�G~�8@<��1ض��U�#K�a�hVK���9G3o��2�b�RW,0�1�B3sd��c$5��Q��@�W�n6�xy]�_��Nox�~d��3w��Ґ��T�����S�>T2#�P6F���{X�B>rH�h{�|����R�R����	8 �]�=k�W�DG#�-�/�>�@OK�E�x^$������I[aw��:�ph�C�	�w���8�Ì��D[���=ȩA����5��[S�2�P�c��-���}bɐ`��dXgSl�5,�aL�+<�(}	a�����x[P���!'��,Ÿ[M?P:��$�-ӂ$s �s���F�(��h'��cƯ�
�mW�= ި�1\�X�?Tk�)JE�u<i���ǌ5_�c9��cհ$��'t�}��>3�"o\TS�^�%�,IR��_�^y����)��s8q��F�/��i1辗:��È"��3[ߛGX�����xU���H������=�=�B�!G�hFҋY�qC�g�j+��S�A�R<C�%6]98�����熘�_�
P�`��o�S�_4;�;N�ũ.?>��-ͷk�����h��Dm��
*���s_����a���:Z:�$Q��Q�����Z�PaDF�>����5`w]0P���XV�U4&���mL.Hx�;~���X\"� bs��>!���a7�1����� E��:�S�6[� �?T�<�����*����[)��#�r��N4���=�D�J����`���4������YY�̡��ry�ķ�&`E>����k��˚���ƿ��I��؟�2��V*���t��Y�i�d��P�b^�L/����'�����f_ʕ���#�弲d�� ���ݪZ���8�_��:i���3F��1�ՙ��z>M񭄢H��L[���+�KoHeQZ�<𓻮x�'O_L%of��N�	n��~[)#��	���Y7
��k���3��T�*��]7����D�*���g��g-?�fl0�<�4�\VF.���]�M��HIp�B�>��Q�m@�'��rgAjd�m��(�,$XW���5C�!�l�>q������2�Ƕ!
��^x��%�?���~��_>�C�����׫������|��|&D��'�j*�e�Le��k��;~��@'�E�0��`�����\�^�1t�_Xaы�@��z�4�Q!��̀��0�ڐ�t:�Q��BE��F���2 �uG|���or%øV����A�5�@��h#LnV��.��1mX��\9K�.Ķ�c:�S?W��TF{
�E�e��O�l.f$�8l��|����"���(u�����l�?���D��Z�3!fݿ�ʘ����H  PR�Q�yώ�N݁7y�2�S��1�ۈ*�"׹��k*]���x�@y�������{��,���]�(r�w����06�>g���F�l�ߎPI����%��(�V�J����$0؜��N�47���Z<ƪ$�f]45d�G���f��sfQ����F�k5ǽ����)��-T��#�5*��7��d�wm�ƗQ׸s��Ŷ��J'�[�A��ɮ�[Wz�\��U���	�Y8f]��"fڲ�#���X���!�2rsZxE��Y�"��"��Iy�Ƃ0oh��Ȧ*柂m�����_K%ړ���!���H��3�}�j�u�o���ző��N�1k����>��Tk��/������M�!�`�ᡎ��!:H�����?.�����=�H��6a{�}� ��O+��̣<�� �#_ͦi�0!
�.<���x�Ʒ�)h/,p%�=��UȜ��]u�c�4����e�����Lu	�||�޿��OӀ���R����&�g�]��o�r4ix��ͥ�{/@Z�5��c����k���g�yz�,���4�plZ7�.aw�>�_ڢ�ɿF��Xmf���(��Y9���n/�l��5�%��ɿ�a�G���)��)�[{}M��M�Dwm7����[�l]LYg
|�{m�|�_7�����BEqv�-��-2���'{���2h�E6І��r��� N���Ǵ���/j�(~]faϭ�
��o<��.���Y���#�Z���͌,1ԑ�V���7�N
D5��F�z��$��L�d�����)��Έ���Ԑ`�lU�F��9���Gzt�\¶��Q�~�akf�U9��b)oKB��>�M��b��-�O{�V����P�%����L�C��c�d����iP:��iC�§��/v�>T���~lk_�����������B�y�衱�y��{e`��k.��=�#�����AN���|C�hL�����W��M�҂��IY��m����#���'OQ_���W���|��'���0��yHN}8I� _ ���J3���͸`�] �����������9��`K	���O��T����M3R���Rٲoǟ�sp+�?28d!$Ӓ�ٝ��(=v��\���~��%�36Ç��Gu�X}�3��7�B:�Z�`H��W�FPiq@�2)Vzi�����>�]v+��3��}oTˮT���4%F���ݧpdn��G���~��X��Q �bMw���
��TLT��}N+�}��VИ���IUv�\���}_F��0�z_W�D��������t�bQ�{	XE��@'-�o\�a�лGy�UJskP����=F�����+�y�#����L�'}�(꩹�Rv��|y���0�0'\.]I%[H\����sD�D_��X�ke��T�I܂�(0E�
,�K��|]fW�A�U)8]���4����^�oQ.)��_3$�E?�7yY !6 Q�  �2x���7\���t�J���hz�jB��\5� �hh�������F��]�2t<��bJ{ߊ��p���Btѹ>\�������̒�|�v�.^7���b0��	����#�s�V��37:/x��$�d�NH���T�@�^�"%U	��X�WK���XcF����$��wDF��#y����Қ�%�ز�I���1C��|hV�h�쫬-���>�tN.��	��G���z�D�ҫ����q�d�]��ޓ�k�[r��B{�t��P$R��W[:NT�d�	b�W�l�N��5���{�a�#�|Ek�D��_]U�n�7�::Nn*E�a��(Tw�9n�H�σ��˿]�1�K��,p�..�ݨ��_;a�`>�k����YS�Hmf�z��V`R��x�L�2�W8ǿ �{aȷP�
Tԙ4ϩ*ϸ����ҽ	LzF	�cs�=8>0����؟�N�Z�ȧ,�Z:�s6��̻Y���I�%�I(�9Q�Y�������[�8~p�Wܓ�Mh�s^�kX�QE��`��z~��w���]u-C|j4ȩ���*��qc��F Ή���p
�.���V��d� /{��Y�f��e�傜����YY9�b&p�-X����fg9��ղ|�S��Q���G���?8������j��~G�b��lw]h�a��A�ä[�׮��z�c�Q���κ�Q�hC�ʗ$,=�sA�+�f�������Ok1I '�݋}�����a�f�B��U�j�6B�����A�X��-OMY4�:��3������;�yٍv�<��KPh��)�
@��(��q_숄��k���mX��ސ��I>]�o4k��4iWK��!j1��U�X;�gL���j���&S'�Ȩ�����-��ʃ���$�����h���3��$�0��e~��
���m�Lt{��;�]�g���4�>���y\Ǟ(�jAb(S쳂�&C�)?[aP'�M2�y�iwV	�5灴��Z\qvG��q��������`o�p�fP��aft�E��s)Ί;bF>c}'�mX��!�Ht3?5��.�x��B����\B�*|Ԕ?zj,e�KH�\�c �
p�GV�{$����c����;����������BuXJU��pi(������b���=I��D�#�{V9�� (f	b�u�s~�O{��/�Ma([�}W��6�g��$w���^����Р5�j�uޥ�Ī݇���sZjIg_�Ѐ��~ebH�<ƛ?��U�]˃{���,���a�/l>�����H��څ����ޚG6��p��#�M>Q���Gv���!5�@�!�Z�m�7ߋ��Y�r��&������z�s.�q;����!�h?O�F����IQ�*��s�h�B�Zm��9��H��4�!��	�L&[}��0y7��}R���ܵT���9�;�Z�K��9O�t�M��{�쳥�(5y��{�@y;��@�f�h�ĩK��`�5W��'䄼�+�G�]����`?%h7x� dN�]ZfKv�Nc��7ukx��m��uU��^X�Uǁ��ȇ*���94A?j���+�+?;m��-<��}v��":�sB~����3`C��"^b&�	6_�\޴�PGzO�@,\wJ�:�,3PN�zZ�DdU-��q�%&�߾:�% �m��|0���QD�ۯ{e>��:��A�/�*�DÊq	k��
w�U�ǝ~����u '��}l?��F�y�Qh���w��(�9�E/&�*:��e���`R������FfB��黙�F�,7�`i�wJ��CC���t57�ӽӼt�\�Up���C[D�J+-$�oA��Z�B��������2�SO5��Rd�Gi�B�y5d��AB��|�5���/������c_�v��z-�y���o����}5�-!�s��������� �ޣ�P��a�+�����ot��k�>ʽ�h��Y�} �WO�*�C}ǖ�rG��_J�Q��6���n6��dH���2���Y���+r�X�+leCW-!VF���F���X�+��]��a �$�D����q����v��*2�Y���M���ҌM5G�����Ի���N�P2�1fIe���q�G,�D���|�ĥ��Gr��k��'�}Qꩀ��m�:�5]]t?Q,�a�4_gCx���wp�mB�5��~\�V*;f;q����PkB����͠��~�^�P9?�2=��+�~�A��tŚ���T�*��x�AI���;����~3�#��*�lҤ6�2����ir�,b�l��aT]A̡��6/�#,/�;���afiV��ˏ�h[��	��_�����uξ'v��<"���&EF`��h�t�X��ȟ4y���գFc����������u\�>r��q���|d6�	�n�Y��L���K+�G-�huU�+���L�䚂F�=`@1y)��}�Ku�N�
�<�$��5��?��q�*A���]	�^w��� )O�(�yVfk6��������;��D^?JCp*ߛg�"�c����*h
�.\EMb�>���."�
�}�v�����ǅ|1�LDf���%�`���~��g����!���O����]#�|���������R�G��,L� ��dCQ� ���-B�?�3�bJ;=E��rȷ5y<��R_��XI�{�ǳ�ɞ�EW-5l�����A?b��+��[:�j~ .s�P�o�v�a��m!�?�\�^/Ᲊ�Lyc��qGD�KЩ垫a{�Q�x�.�i�1����+���
���<��~���'�'��\N�Ʌ�]���u�����۽6}�3�=��U! ���﬜a���A�t5��{�m��l;y)u3S�RL �lYl�R�F���*=E���>��X�*���^��K�q�b��#(0:'�He��7�J2��eUWaom�FH�m�nܲ$o'��{�1HS�D\�h����3�!Ĺ� �Ѕ��٫P�!� l�ʢc�������g�0�Pz���5dm>���NF�j�!4W��Y�g��3[AP��G���P���a���_���}c��4Q	q.Kjd�C����G0�*�ֆ5�|$:�[��k�t��*<?b�>�֋3����"u�Y:V��!0����=��1���~8��Yf�� HC�����]�BT,��yG�p���"��x���7�W�(#t���݁#P�����(Ё��
��7��y�i���W��A��029��"�N]��L�d���e,�e��T�����~�;���������b(ޓ�
�f�Y�F�0��n�I��xEA��?|�Ȥ�E��>5(�k���[xiDJ֛�y��r^�J��f�˚�ԑ`����/���&1cv���=	��T����~Mr�_�"��7U����Ǎ�[S���kå4f,BZ�s⇛j���?�Lص��ۦ����>�v��f�bI��f�o����<!��F�i�zL���3�c"b�LH/a������u��Ь�n^�+z�Q	��w�	�X����u�5����,�O�#���knU}��sR���� ���h�T�&ybm/BMJ�r-�V���'#H���9*�X~�(�|Zjp�6na���� Q�n�)��"�j9%���~k+y>W�H
���)�5,We���'�eq�9�����8EV���c�\32
6*�FҞ;��C���;�L�����R�w_%�%�qy}�v��?�)4��(�"�WB�
�S=���;B*�fe��Ǣ��q�F �����y�f�4���x���$�M�o��.�@R��#���IRV��3պj��0�7YC���p���`�/=��	�#���PFy��_7،�N4zg�X�2���}j����nm�'��d�-���g� ��z�y�$�m^h�Ӯg�&�8�zW-�sy�D�[���ﰯ�ӍlѲY��k�?z�MC���͈䛐�d��gs^���URG���S̢�*������U��q~���-�=�<��\�"�@�rnl���:�q�� �T��N@Y�ƣ��5V<��O�&ł�yJ�6��f��Y(�2ǳl�F03k��2���.�5F��<��Ai��J��;��ÅRQ�3e�t��<j�F	�%�
ɢN�Eʬ�S��ٛ�wD:�]c�n��R��K\#�a�AA�
�g�;�n�|lG7���|N�˩ 9���!}�Z�@�?�,k[��i���	�� N��`}��5Oh��Z5�r�"�+L��|t���A\٩�#��=b�y�@Za�"�JG�Q��J�O��g#�z64�`b�מ+e��Rp$ɸVձ�_��1��E��
���T�jKf�Rz�Gݙޫ��
�!g��^�� :d��8�S�0J���ѻ�eԕ���;x~�Lb�%��Zv�Ղ2�!޶�r߾��R�y����0����S������s�*��Nt��Fô ��0����I�d
!�Af���J�p����w�}De��u� �>�B��n���C���rj��0P����u���~	�V�i�� wvT���'��D8�a�i[��Z��2�f��د�,�]��J��h}����i�=���k�4�u��^zIJc	-�ۧ?���Je��� ��?��u,6��/���p��k�䨨��9��_�0lR�T."���wy)T D����ًxC�#����^c6�F��5�wh80ŋ�(gm�&�6ܡ֌�F��O��i�+�Fu�|��c_Y�.�?j���W e_G���U��%��0U�������'�=��Q!��:��0к/p����h`�<)H�t�Ó��o���8^�=�ZԚ�6�w>j"���;`��%'�MjBSP;����G]Ea't��"X�U@a���Ӫ�C"�RrD�q��U@�:���~j_2/ $ ƥ��c4ߗ�yo����y
f�R~O:_�]�5TK��<˰4i�c���&,)n�f����m��~�ߜq�us:�z\�Q�Z)��t߻s
��`����fڂ� ��4|�8�㑵;�T%P�G§=d�00�����i��[���=��u͋��Au��� ��½�^Y{[��Ǧ�}�K���]�����6&�m��jI(U ��#~"�O�h��o���?E�o(ik���e]f8�*"'�2���q͸���m@�L�8q��`�#��XB����'R�K��h����q��Gػ^���	r�tU��[t���В=y��'G���y� �����u�R:9��u__-�r14_@�w�0;�v,{�� ��W�'�����g�r�7�T���,�-ͷ�YZ���k���m���ө>7jB����5[9]C���I~���ݡ��#�{��n�e��w���8��I_���c9�^ze��"3b�Fo��X���Ы�Ko�[�>��l���Ag��z�}揺�o	����̓z���J�<L0�agC�h����1{�AN��A�~��g�y��E���e�C޿�� >�Hn3�WE^��d����i6ŗ�<��/��Bе�А��4�̤��]m�M���X�. +t`��y�Qa՛ԏ�~� Fn?<i�2��#���������\{$�lc �Yd�Ճ^`@aq�����p�.k5��?]���ޯ9�Zq4'"�KC,���L����Hw+�Qz걐�L!��OŰ�V�Pnv�sO���ZS�T*9�^s�Ї�Z�K5l\�~\C�� �4|�������(:�p�o����po .z����	B3��6G*w����oʬ��)=��r�Q�~�� BG$:J�a������п�t��l����˵�[����Ea���Y��-
��+1�r;��m�@N�8Si�_c�Aƃ�Q�(CMq�4":��z�#��2��ǩ�����#�0Z�eK�M�.�09$i���|6�ǯ*veVա��O�$r2��r�G2O���t�?T����k�lcbD�. y{	`�p���w���ۿ �,_�L�7���x&�v�e�ʷ���z���L�~��Tg}�pp�c+�P�D<Ŗ*�!�O��$�fg=Ůq� �$d�-�L�UP�ap3l�1y0��R��pBduv$)���5�C��i�/L�`��)UَZ#��_����j3ñ�",��|�W���`t0��]u���)�g��N `�\|T-G
���P�����cu�cjl��|���m��&һ}�0/R���:�M�|�\�]�����z��%@xw��f�i��t�aq����=}Q7p?������_����y ��jȯ���l��v5���5��sKbb!���a&���L��0���-�u�BX�I0��G�"�/	0G��H�(~��z�/��^׈��H|�`�2&��-D��<���c���KHBE�>�i|�r磛k�D�����,~s�
JOBE�`�lա��ѩj���*�r�?������;���3yc	2e9��A�lLZ��1���L$��")�Bc�o69��~v���hU��yYm����� ���pEg�Oa{Db��	D]+�&a�"�p�Cα����GJ�߁��.T��<����Ț�n��SͱO�V#�(q_�{�u'b��߲��AN�p׿'�:D%��G�f ? nM��R{sd�&�J�s@I��5���k��`�q�L|�pn�Pk�Q%�eY>��0L	��X�~��:���{�E�B�K�lt���s{|�r��<C�j��� $�)ʁ):�U�~{+!zb�`�r���@���{��A���+�V*�@��ܟ����>�}qZ��F�R�|
�f��j����a��{�Re��5�6�LE����|�E�a�Ǌ�w����'}��D��~Z��4�=n�x��.�о��{ˀ	�}�ђ<�<��m��\��l���S�	L c�*[�������: t�7K)g�H���F��Q��A��h��Did���Ah� ��@g�F�DѸ�5uJ�N/9Ы��Y����FO�#7�#���<5�����wf�O0�9�2������}��iԂ�f�r��2-��j�ɣv�}�x��;�"l�R3���V�r����/��6"@����G˯n��%+�j�&�x��W�-u1��x[�]Wyx��@�Ia�iP�Y���>����������j⟬*ƚ�9�s{���D�g�u^hĴAUh��t��dj��&�����`��;��t]it�������FP�pfmy�~Њ� ���J|	e<X<;��F����֕@Y�y�F��r���hϲK܍�A�݁�N�\g�H���S[�2�� ���&��@����e`�������� oy��AC������"B��*�_+>Jq��_=��u��l��sGBZwT��%8k�X/��RSznа�������0�KAT�S&�xtw4�A���;��������}����1��o��Ε:���S��i�����a�c	����0�8�9(���R`�,��z5H��W���պ�p]������5�Q�߲A �K�F�[��t�Z��%T���JU��~'�n��Nz���h�@Q*<;A���B�U��
�ː��e��{!�*����N`�U^Z-xܡ9\�jr|D�2	��$[���@��{p�KC����2z3��ظ��<=�*�u��a���X^�OE�����ᣅ�ː�ǟ�~�H覙��s�2�-)���YN�������9�o��B�!M��{��W���{�5�9����Q�/��M=���N�o!fJ�#r��Q�IAAD&i��R��Qi_ ���<��)g���r���㹱�.A��3��k�� ��kW���6v�-] ؚ<���}�W^hI�+֧����]�d�����
n��G'1HQ�i�*0Ob�I�ӡ���@7���{�%�O�\@1��2=fF8�&��d����}�E왜�jL������#~�oߟBd�w��G^MB�n�(��5�J1���HL-���EqA�B��I^���K�{�$ʤ�(Y�ğ���n�e���8ㆬ
�Q"Y��������^ڃڊV��Z�����^(���i����Z���=ג��2�����
�#��H\���_��d�T40�C�	��V�%!8gD���5~koY����$��ˀ�e��e�y-��Eh��y(��!ɮ�a}5{6'5*n8�M\���Sޛ���I@��;�NZi3	��[���:�Rשչ+��t]R~y�L�3X�͉���0?I��X���;��%L6�zo��F����y<r����2��3�|������j�*w����c��B6����$�4�eu��Ũ��!A�x��9'��GUN��m��_XK�-ޜ62IЋY�-s-�{{�.Q�H��:�0	���O�\_��M�l'?�V1pe��;G.U����l����v J���R_���!��k��Y�ި޶pQ詩:߷��1/��	t�4�Iw��:f���{�^��m3��hS_���-���*���Hp03�X͓�:�C�w��;���N�x�B���xa�������vVӪ�����_r�\Tg��Դ�,f���V��/�۵�M�n�x79g"xpk���[DB�Ϯ[�������:��~wD|���ծ�ׂKg��)E�=�_7����sԳ�H�����8�o�@Ѫ|vb�S�Y�i����,����<�ÇǢ���Y�'�.q�ah�9Y^E�!���>���{5vغ�]���ͬ�}�k�=/M��Ň�g��x,7,&k���&̮(��zk�R��n���sU��ͳe.o���<���	�~��⪗�i����,f�����v�L�	��#���<+���H���\sf���X4��KG��	C
�/U��o9�г��e;�%�����1AucC��3���/z�)4%�-a�M)˔?�� Rm����血q��fy��[��J���۟f�P��Z`mZ�8Y.t��vc_��Ib_�R]gɭ-yC]ͽ�Gڊ�����s*�_��KXaM���k�L�ه��6Q��ܬ���NRae�C�Pu?�8�#o��d��ϼ�ڂ��˭�Ƽ�Vd0��w�|�P�d��Z�L`�U^�r�i�X��	�S��~ARy��I�ƍ���J�ک>�s�H!h��kƹ��{UIj_��>T�g@z�Q��G�rN�Io[���r}#����z�����J�^uO�'�*G��GW�f�{Ͳu�U�����b�����e�GQ2�=��.>��:J� �x�H�����wF>!�Yv%�Yp�uH8����/��=��9��K��-U�ٿ}�w´�vbX� �O�����q.�o�v��W�o_��mN�Ζ�t�ԄT !űܓJg�W�+���F)u0��S���L��\���{�H�����=�oMc'��4�N�����	!C;B�t��R��t�HncM���,�����7as�b_�J���l�J�����	@����.�	�3��d#��C��[ZOD��6�$�f� qЋ%7T�r�D�[~7�����^฀�L�Jy���b6V�5��`�w�w����Z�I,��⣀X�G2O	"�J��L�J�t�8J� "!��������������:��`U�Y�D7J�����ݿ5��KUWI�̱Q���sU_�1P��0wK�!���=���e��C��m>u�D�J�����^�Ϣ�|a-�������ؤ�U��ٳ��"��[c�8�r�C�]U�
�z̬>a��o����Ć�cy�g?�kr�r��'��~��p� ��b�����-���8Y��;������-l�L�wS/q�>}^� v���� \1@�czο'%�ױ�����P�-{���qA9HާR�DN�g���OY�1u��o�9?&�a���П<j�@�rk_KWYj~/��_��;t��*�)��7�'"'������6�ߚ�5�v��Pzk���L�ɭQ�B�4�.6L�w�4?��~~������Z����g��+h�5I�=jn���(�֎�����6���'�O�>�T��3y)[m	K��;ԕe��f�&����Cs��b'k�^8����N��S(�,t���p*�c�w�n�)� ��I*�kO�����'1?2_��p���c@=���~����P���h]�z��7k̕��,��AP`y�S��z�\�u@T�n�/!
�&�ylXW�4�
](O��k+���G=/hv�BBkX,
MJ�Y�^��%��9���6�|�fN+���u�� ��|f�U]���o'F���B[��Sz�Ϭ���z��N�����s7H<Y�s����@>��B�/Q�:M8l ������7Z/��F,�����V��#�3�%���3��h ���^Dܤ����Z�~��I�hP2$WV�����Љ$�~�֡��ّ��cl�ky��@}|�V�=�/�U2u]���>�"(S��56�ڧ�͗ҶU��S_�a�SR�|4_���D��Wm@g��Q���AD)����!Dk�k1�����gD>��ń jWN�����iG���8+q� �De�*���y�� #�!H��+����-KjV�d���r*�X1������Ԣ$V��L�|��qNeV9���2|�z|���HU�-�<䀛�g%�zQ}����dTd��;.+e2��Ig���;�Q��l�)L[4��ۑ��*��~�A �<5��*�0m���-�N����%�ԣ�|�s����w�^Yn�\x���;� ��,��'����n�G�x�aƧ�g�r*��A�1��;�Eԏt�������)�"N���%\�B<}�\oyo^~��ڸPg&ǋ*�jb|�N���R�����A� TZ��a⊭���ۮ[;���D�U�S�-��+��uET(~v��t��-�x�l��kؽ����&��N���<@J�4Y ��?�	Z#u~U�O��k2�)����7<S���k׈�KIquȧ>�if�{�b�%A�N<%=�ґբ��<]���} G��E3�P�Ͼ,x����:]�W���?��h*�w���K�Ebm��arx�>}A݇��u|��A��4�ؾ�Fr���{c���cv�(<���K;O�_vy[�g�F*S�:��nJ8��
W;qN����5m��������j���@+�.[o����z�)���p�G�2���3L��]]B���;^�������P�q���"$�w�"co��0�~P���! 잳�l���7�>���%�pu��}���׹88x&��t��P�� P��q���,�����^���	J��A�i�נ���s�i����E�j�55���[D�^!��MA�sȻ��Aد�ә��;���f��1���_*r#�s�Ҍ��l��i�@�*r��{ԴM�	\�3��dOผ�� �v�i�GV�Z46D�:n�ZLs��Q1H���V��c��y�a%����/��᠑Չ�Ԛ���b����W�(?�z��R�e$�^Ǻ�@ft��Es:�B�!h�!&�{:��Y�V��n���a��!�;t}����5�������Rj���� 8��
��i����M�����S�U����@@���[w�uj��&W��u���E{��~p�n�`�������:��ײiϪ�� r
eIEb���y��: r��{�E���82sE0��8&@�J��(H�aT@��@���q�$ �b���t�A����6�dhr��9U����_��/��Z�.ƪ:g�����g�*��16��#�>B�ƭ4O](�D��y*�W�s�Q��Es鄉�:W�?Ij�W����������l|��#OU䢸���� 5N�Ӥ��Mx�!M n
����/&&>U�F?�Y�8�>�	��5>�Hf��v-t���Cv��u�Dɳ���>z���'z������L�Q
�D.��j������M��hc�����%PN�1��I>���^�׊q+O����!��|��Z��dX4����� �Z����(�N��ڬQ�����vv�	�j�A�ϡ�fU���eUA�~''oA�.�$u�fs�ʇ�R^/-F>�����Z���A_Y8C{F��~0���.�^X���@R�Hq��H�C��&��7�[����(˗�i��� �j�?P)��ZCQƞ��4�F"�͌��)��1�_R�ߢ9/��ާj��C���e�Å8&�������G95@� B�I�8��4Lw��|� ߆�K{}!��c/���A��-���N˧�xl�|>e���U�둺@���	����.\8���֧�t�g��`��kLl|��8���A�����&�Z�m��q�#7��E�86�н�����PY����>:o� V|�&��1�c[�����|�mBڗX��:m}yױ��HȒ=� Ś�q�}Q��uh�x�xg5tv�Ә�9/���ve��VQ$&n���8�X�n�?���qA�6�+(7��6���2�Kq\:L��1�����tn��.�$G�����{��)�/���F�MT�-�����E�s���pB�^y�,}
�g�o�̺,|������X�N�;����]�ƛ�HJ�7�ThtMAr�n/���j~�~4����P(����(�t�p%r�vH�@>��~���j���Z�=���:�͔�A�r8�H�@�M�����9t��������?A:o��)��ǫ����zty�u"ȴ����)k)c�S=�HsG����U�Li�N�����Ȭ�e�B�dz��5���ª�w��ɚv7P*��G'-�*�� ٧����n��c��oe������4��+��<���s��*�lu�	M.u7K
�zϹ��k�d��x+I�.���bD ����&�Џs�0e�u��N���}�KA$s�x�	s �v�k�(��d4�&sG��u6/>q?n���:��v�>0��� �����Xؗ�M��~̧�k�ae�b# ��_�����P^2�R�h"��l���S�ڦ+�=�O��}m���?N� �-�vay�*�����-yF���!|��#Ӑ�_�����<NG}���AX����9����C�&A� �Wޟ�(��:7ydw`�Q���RՕ�gzz�\}�|iq� �����$��@z��\�r�U�#ਝ�o�������vY�G�~R���@i��;s�별��8��Ey�]����/V�|o��]�$�����+®~㠲6�j�w)����{ޔ(#�0��s����d�����j��|��N�/�nϋ�W��ԓ&��j��WN�� �Y��Křƛ ���jεq����	�╫�"h���%,(=�0iw�Ջ�H�w��#�������p�����g���C�U�]�ۖ��{�QU�j}=�r D����Y6�9է�Sչ��%_J��̏ �	�%�,x(����[H:ICtS�&��.�y�[��s��_�207��W��S��f�Hbu�.�OD��Cn�#�* �����^���R��Rl^�U��$�P�{.i���W�#
R����1UP*�<K�{46Jy-{�����"�����zQ�~k^��O�Q"MZ؁� 5������;���:*(/��C��k��(Q�g����MoJ}gG���S�}%L����& h��AR_���6�__�vr�RP*,n;�s�O��MM��9s�> �ȇ��������W}d,"�#��Tlr��]�ڰȿ �ʾ�N��.�e��N�$�?B�?zT%[P���T{��K,�7;~K���q��-�������������'���ؓ�ҷl�������h������cN;NןY���iX,��o���^�s�JYӣ���f��n$q�Qy_%�ڽ�t(jjEU�%o��u�m8��\]�4�ƍIe�76_�n��6Vx��Im��9|�[�b��3�S�[��W�,��p����A$Ҥy�Ło���K��`�X _L�rX���t�h1�����7�8Y]���&�~>�섋'B�]�k�Ȥ�Ak�M��i*H(B��*�1�e�!I��7���bV?�Oۓ6�^h�uF{Bq����	�U�N E����N��)p�6]�����n>�E'�8��S���!���>���۞[��I��EWE�"��Yx��Nۮ�>d�9FuG�ĵ��"���yu��K<4<��%���g�K����V�Y��S��J?��lEsI��v���'uS���Y���Vm�G򷄽�sm>[@9���ѓ�9|���GWzT��)�85S�͈l���D�����:��,�r��'��%hv~�n�Y��4l���Nhp���\�l�Y�� �'� _8�#'�Z�/�#���ا��9��[�p�E��v/FG�7��>fe˕\OJ���ߟG�xNMJ��e%1ڃ`'R&.�S�`�B��.�Q������-?���i�w�oD���?@
�0�x>ٙ5ݏ4�(o�m�{MB<�:�v�{�κ	��V��Y)��k<����n��o�^�K�B$���&QFs�u7��i.����ȁ��吢�6�!��$6j�i��،QX�X<:�� ����y��l�~��gAα��!�-��_����z+l��m �B�?B�*��Mg�n�:ru�˄��n��]�>^	N�>�f�����+��uҙ8_�''�zW����&�]l���nu��Ǔp����;�ޭ�F�|ҝ�wϪ��/�m���C��L���7���Y)s���'�YI�E���0������l|�!2��:���?{��q��sk�r($�ԇ��48�~uJѕ��#�p~��T�C��l��;͢���z!6^G��9��҇�:���u^H'I�H滤�J��s����$7.x�:?���kI���y%�9Зڱ6zQhf7�.���L��F/���/`FjQo����&�Dy[�f�_I�O�)�]ob��߀����F�6N���]o+7{�������,���g32���e���/f2�"$12���yO���=	�p���U�Z�riv8=���2i�2-��[$~�߱���]��p��BFQ��rH� S̦ӓ���	GA��壟�k���d��- rg�p`WZ�DMsE�#�*����f�e�ꕽ
ܥWƱd�T���)1�(����7T$L�����Nn���|d_��z��z�����v���q�1��NQz��B���k�B��]���G6�8��C�J�A�{I�y=`k�S�A��B� ��w�]�?��/��0Eo��>��e��0��c���Ŕ: �;+��$��o������O4E�먼=O�6mH��<��%������%+���0@_M�	'��M�;��?�I��p�$ǧ6�F�	� i�]Œ��UQj8G��с��y@�#֖V�����z4�P�y
t�g@���q���!�+�S�N��y���SB�̂i����]��2�W&��خ��u{%o��x����;E��ԣ���R�O���J|[�@��P���Y�q�Z��-��d�C�ss�u�-�Ps�L��.A�Z8\��g��Kb-�^fj3�,�31��L3��bq�z5�_q>�t'��3 ������,X�@&[�Y}�^�Z���.�7*ڡ�aa٘?��&��UVeFa�T�.Hfm5W2oI�����3'#�_��LB�\�d��rҭy�6�4��{pN��C���{d�_�G`H�X~m_&A���2Ǖ�fq�3)���,�/��.�u��	����.]��ܩ��+�u��՟Q�˷T|Q*��`��(�&�������(����`���9��{�F����Z��X��<�����=���R �u������y�*��:$)	�o�Q�R	�U�����he*\����>�Q���c;E(ݥ$�4)�q�{L!gŁ�͛	�E�w��D83x����h,,��/i:�A�@�w"�]�u]�ׅ���63����|ݾG�,������欌����B�A�]���i奡��^�A_������3���ѫe�7��<(@����	�9�Q@�M"F��܀[*=F]J՟���I��׮a�1N�%-:��T�䖿p@�#6�v�~z��0P���߯��G��f��~�"e0�qFSO�0�Pl��ˤ�Ԫ��`$�� �J��S?􍣀�$W��W���T:?O�É[Օ��D���m�!}�-��ֿ�[��B��2#�9��>�g� �n.p�(g��<�'����B���0o�%K[��a^��2�Sv[���a���[ ���Y��ֳҗ���MuB{�Sq.y�Z�' ������:���Z��J<§+O�AUZ����Q8i͌����'p�wO�_���~,3�N����@��a��%$��/�vP��[��u+O��i
=��r��ڧ���D�r�mA��#�-�B���d-���*��S� ������,�2���L�7�%�����S̩���C�N Q{!�̯���T�e��7�~�N��p]�ج%E��I�pڀ�jG2�����*$��]I ��$��E v1u�<®��;�\_�E2lC
��vg��\C��K�;o#pY��g����g�k�J��9X�j3��� E�\w���g�*�z]8$��"�bg ��o$)�Lʐ���}�AI<�i
w�$>Y�ʰ��}� ��:��?:|�=�ϝIN�ݏ�D��v]k&A�d8E>�����|I�͋��K<h�v.:�muf%�:�58�ȧY��b�6Ԁ+<du[�x�q2��!��[W��iB�<�� �iݮg�����ӂm��� wn���ɬ%�\D9��-_]O���h�uM�b��� /��Q���_F�$�!.�jZm���w����_qu�K�ɡI
����	�=��,��Q�v���p!��,����"NN�~ѵ<d� ��RAx���=�����k]�ɇ��tt�
+�뷸�;�S=8�L��@n����T���֋��R9�u�#(��M��j���T#� 	^�Oߡ݊�C�=�i#�����#Pa� G,!��}��7��~*���������>�-�b ��:���.j��FeoWQ�j�-��e�"[n�-���Rn:0�Ӎ�^�$B��^�(���6$ܧ�V� ���q�t��b�U�����pokK9@�:*�j�������Vh5���Ay��)��n3�X��^�iZ
7p�J�ƚ\P�A��jƢ�oc��c(���6��9���ihX�V9�|c> �M�z��3e����+��8��Bn#�w&p�����Z�d�yU��,������a�'m&���~4x�RO--�+�N�3�N����E�D�"��j+�D����j\�Bg0l�=5�(g4�ts��+�>��2�Ek[�	�v�ӕ�od�*�L/��i��&�/�f��;�p��$�f���j%�9��
"`�2�duzm�()m%q�4�irr��0lX��{8&��৵@�������ڳn�l�2�����+WϾ��d}S��[BK?��o����Jl��$f)J����嵻{��C1�K+�*3�cZBJ����@�ì�<���89��]C�&]w�4��Z͌��\���cR����E�~f�0���U
�������BPS(�cRj����-/�dBAQ[~���A.���4��*0� b���w��0��n)�_��K��nvjN��%�҆k�>
~��>7k�S����~q=��V4�Ք�;<�����ͼ�f��#��t�#�eU�����g<�T��B3��Lj����aM�' ��6��k����/��o������ �Uc����r>	��P,~�罤�$����G�m�r��
d�$�/I�>�=�����B6�0R)~�����(�ˋ�l�S🖟kY0**hU�
X�%��e�R�(�K�j�>�,ml�P(����8p���4$r���mEd���x캤�Jc�1M?{.�VS�8�(��+ �Ճ�����6Ȋ��K�.G��}��\�|������uP�(Gw����?�v��l�X�ȧPTV���sf�	7Ɉ#z�nŗ���C��n&��ОH$w�]~���P�Dyt�w�C����g�3��t��>f$T3k�9�A��9�<8!R�R�gpf��:��Lu��F��:D���+�����u�����W�&�1&���6C�)6���c�DT	w�By��8�����~Z�z�!&��%#�]���$P��w���ؿ�I��/�� ř9�A���֬��%�Z�{PJ�RJ*�m���*e;*5� 
��U|��P���\�&o$���<��a't'��.׿�����vγ|�p��ˏ][��>n���FҒ�2�z8���_s&6Qޖ���w�we�5���u�"�v4��Ш�Q	��T�v�����p�'�]5i
���q,;S��e����dD��Zy/�6%2!���˼�|o ��:y~$UG�Lo�7�[w(A�	[��ʙ�	�A�dX	�7o�dOqԨa�+����#_��d0��[]�KNÎ	�&�8�39���}�gl2��|���|GM��Ʒ�*�=b���˾���^�%��޺lo{#/�-�$O�2��Q��݆ks<
*D�^�~�O��T&��8ny��c=t���Lv��QH�^�U�f����w%<���<��δZ���<o��w�.��!)ÉR2��B\���݇�SsAƾmf�Hې��~��Oq` �ѯ�ߟ�;�x�!]x�	79\�������d�Ƶ[�Hg���s\��:M��D��g�R�<y#�㰠(|I�e�,m���b]�T�	ŵ��2��.�}�QA2;<�n���_�Ar@u�9��Eƪ-��7��7��Ѱ����%ʿ�i��DK�l*MH�i���"�k�9V~�
;�3B�o���ʖ~��L0��$��L�]sȊqa�/?@&�؜�ޚ�9< �N���GM�7�n��b�$Z�� �4�Sϟ�愘(��*X��aO��?r�PK�EFTJ��������!��O `��
O�qUd�ۍ�W�5�9]�b�LR��G�	ܛ��Q���!h��o,�|-ކ?��@|���5��[E���a�v1���Q��*ʅ�-rی�KC=���@���F,mzE٨xA��ī|���p*�F��6P}㇗�P�_\1���������N$�k�B'���a"w!+�k7o�8T�P���V~7�:�i�U������ЉUO�p�8������t`�o�Í/I�+p[z�C���7���'@��`���cΗ���3Q���D�(�*1ݺ7?"��[���O��p7��U��H��#/Hp ����3�q�<D�|B������w䳦F|U=Yg����̚�\iN)-�b߳dt�4?",~�	x�f��g^t\z<���-��~
�]��vF1�&�B^�|�_����"}��(Jf�qqwo�6��j�,�qH����'��I�.~�-�= �~����Ȧ��D�W�#.0�w;���Ӌ�07q����������)w6�־��($�M�������Y!̰3]H`��R��0�;!՘�N� -��;�LC�i��g��_�Na�2=rF����m���-<�&5�2*D���������;o?L7S�F����p�F~�0Ʌ������h���&��#�!�թ�M�_�o�����1
t�9�,��=R����_�+àl�]P����{שZ��H(e�ȘC�x$�������M�����<� �^��J��_6_j���.b�Q#���۴�y !E<��<Cf���#��{�<�E�p�����ʰf< ͊�˜/�S��HNS�1*�P����R���������d;7D�~�Hƒ�9) �w@��[8��ҧ����r��Mya�nٔ��i]�Br,�'8�<�y�ϓ�֔�;����j���V���`?#9C�ÓmV?�@QA4J�n��	n��Gc�.aw��,D�إn���n���Ƀ�=IW�P
��?�b�$�l`�W�D(g�����E{�p����s�Cۆ�|n��,���e��tDqq G���[��=�0S�뛋b
�y���m(w��R��iE]��|9�i�9�j�:Y��3��Q,If]�t�%�q��T��Ɂ�46�w{��mvK��0��5�0e��:��(�c�f�����Q�$�.�2��E�#�rm&� )+�\]���߿ϴ�W�A�`����*�����^���2ZO3�>h�U��K�������K΢
�T6A#��8�.>�S>�9�ӧ����B	SW���aH*�V@��N�t���X��&�����Cn���{j�C� ����zv����)_m�����n7X�k�3᝻�����L�y�8*8j�x�DW���E�����y�na5*���2�y2�ij���_�f���c�qt���I��6���f���S �Ct���H	f��m��δ��7`%#�e��־��Y���5J奾���)���}�c~�!`�	5N�������EƢ��?��d-�c��OTHUeW��G`���Y�� ���Rq2��<��\���
K��!�֎��i_L�Fk����Rb�|f0�?G$�����ל����E%��@M�$7֕(g 翲��^�G�d�~��BsBWT�H*XB��ڭ̕h��f�5z5% 
� ���7(��zRr� ͅ�v^5A�]=`��� !�grA<�!�'����im d ���@v/�ε!�kg��ȡ�������3H8d��O��ѵ�(	��4�D�s.b�M��
�D�l���,��C�zγ	�����郞'+�	�fL�}s���*�����}p��?,�&����T�w��f1�N n9�:8�N�?w	0�\��W�
P���Eg��@ß��m����Ⅸ9�~,|�+*I�T0Cҁ�<@�Z�����G��a?��fDٯ���ֺ�=��2$�"�$�L�h3Y&��O1j)�{���ֿ/{�!G����1���m2�.�����o�#԰]$ې��/�C��F��{r݌	T�͉W!ַ�'��)��A�1��5l���x�U�L���fp��-/��4�@m��6���܃�2�����'|�x��nm�6�~
S�轗�s�K�@6�lLu�ԏ#�9�  b�yzm	Pa��b�� h��'w�Hf-+I��j>�7�6��R0�T���œE��-BD-9ņ�5*�`-dVW���P3[+}�F-#1�M
@/=є� 6�B�_z\�{'��`�������j�:#`X�d`�%*E�	^�z�)JZ8�
 ��C|�w��fd�G3��R-�� ٽLȗ�	ڇ�����N�:���*d�h�^דe�"_���icV���`�ȔKX����"����(�h�Q�"��xBsY�\��P�~dw�^e��|�SE����,S�n^:����3mm��$+���vzX�E���F�Ov X8�ι ���45��O�e��õ�d3�G(�C�I�:c��m֮!�P��\��5j��M����}��o�=��
d=�9FC���"�]��)�#`B���O���,�8�z�;���;�ȁl�q��D�̲|����[�A ��������:>�������c��JK+Z���� 0�-���Y���Ϭ,� ����,�}�\����}� )֞�}�����������
P.Cy�W�K��k��,��v;Dz��M5��w����E,�"����f�S�|�" ��?���j���w  ,Ew�pml�`~C�]���Ba�L���z˷�g��7R��o���k�t�e�e��ۃ�'�1�o3A�� �H֝�����"��7,��n�[Ѵ=�I�E͙
�"�{U��k��]sr�qS^`�~�r:�>U~��o>iV�Di�+	���LO<���4loe��=�hL�9C���ٞ �\u���?����@��!(���DKuI!���򲪢���@V����Ϳ�௷�� ��w�&�G
GQ]�o��L�{��|�����^w�j�N��[W������bs�"��`^ 5���k�Ji�Z�h� F�?nY7�_�F����ЮV�@���-W@�;Fq��;ia��~j�ϯ4��v �f��jAR���/��a}A(�Q��&���!��|�u�M�
>6{��m5|�du�pd����
1��] ��A���鐏�7���n/lt���|}<�7��O�|�Ŵe(��\���@.�H�Ȕ�L�Yl#q(�.����m�@�Z�2�i�:2j�ζ�>�fBy>#�X����}fT�p��Iv!�Wˇ8�OUz� .��u���$�a��Iݗ�Y������~|� ��oi��fQɧz�Wm��X{U���?������XW-�����^ܳ>�b����=���y@�Mm�	j�i`{)�olEr1���&7/�6��*�2���+�w��}|�Z���@�w��I���F���[�ea%5����pdgi(硐�ζ�F^p�һ H����������O'< \�U�� 1��`�0���#�O���?��Nb�1=0��Uo�E���i#����b�"L*:}q�����`��6�г����8�{|�hw❴��1�8��\A�Z����#��K%MjFAq�L]&C{�}�$�F`8�埳��R�vf���Y��UJ��!s ���p�z��8�1(�E��D�,� </n86�t5�H�~�pfN�|�q/fk(kSdޅ��P�a%��?�e��qf��)D�.��<Q�X>h�X>&c=ٸ��X{:H8/����㏸HKב������������xwD�G �{ԗ3F��ڏ�o�3Kb��o��K�H
�Vב-��K�,����Pi�A&�b��÷��Ϗu<K_�K�q̺��S�l�޻�9OՈ���������4�u���颌��V�x�\`��Hz�wF��uO�������؟�[�d���i4�/>6�惘�Qr��pȪ��r�kౡ�(��kgb���}h'�ߊw��/�M5�h�ixAw]I�u9�Zҝm����D�%ŭo\)S����K���?�t��	����˭��-\Y��9�t���<㿲
+��+n�=o}������er�Y(�T��moV�)��ɠ>4z�]�Ԫ=�H�P1����y,>���n���(��+���x;�Bn5 �*rn�
Z��+u��_`d"�'�,s��C�(���5�~�ɣ����Nem�W�����5m<G���TI�x��=���	تwe�Vp�;S>�֢� +��n�Jp�a<��1�v���0���oN/x���@D;.��8Ca�|ES :eߑ�f�?���(�_zI�Ɇth$Å��t�k2*d�Ζ���'��]Vti��x�G��f��|(qu2�7!LN�cmlhq�,#H^�b�����B��C�48q;���^Fc[��
������ן���&{]5X�O��V9��ڏQ+^7{�J���=%
K�M�x�w۸�x�p��@�o.����4�b �DT�-�'Ʋ�M[�<�u<��dp�PEc�2�%����-�(��������s�{p�����[ ����yY�"�8ye�N����^_���ɻyfI|1 N���7��7��ί4/��0N��p�����~��{}���h�i���Ӱ�k�|L�d��;�F!P�uߋ�p-����zCgI��q[������`y��ȹ�+�3��3���t7���.{��6��
�w��xq��J`V�
h\O��t�ֹ�0��S��]�Xb|��Xߵ��ɼJ*���n7J��3���QI����ڱ���ޜ������?��W����^�yt�=���ª����ǲ�����<�M}!A���#Ul�+��^Ge3��{1�� ��0�g��_�8�0X��?��Զ�bm���	!J�9h]=�����k��&?��O�d, ���1� ���6��a6L���?�o=U��2nl2�pP��h�x2��Gb$|��/��D�y�I�!#"1,��7H���9�T��H�A�j �;ί�6��v�>M�������j����c�$����g��4����-��x/H��O����"Dʥ�t@��q0D��5��?}������c~����#_�)QG���9q�}�9��·���ќ��z��p�!F��j���i+�z8������S-�	t�{K�a�3�YG����x@��n�+�#���A��X �?C7�pZ��S$	pySC�|%�+�� ^��?��Z�8\?LAG�~�a�!���k��������y��x��+߀O(��s2�����u��o\h��0@�2b�ۙ\������x��9dq �"ұ�x<��5+�NV��	�v�9lNSX�� �@7ކ�S�>��4!���7; �Q��dV�F���y��c5��d�<
�o)�c�!5}ݡ��,��8ׄ�_J�$�5�y����\��)O0Q��↤b�~K�����N^pm���VT1B1��!�@�R�_��2B	�e}��T��1/����8Ǯ����r\��(+ �5((�I�4�n����i{R���Ձ�ޚ%� ���*���~t�	�t� �sdj@1�x�'#���R��c%�_���梻��̀v6��Dy\�����3mm��u�"y�m2��?)�f].y0�Q a�8�j���y��ZӠg�=<U�փ�jc$SS�=��A�ǁ���i<�i�W�2��] n��ټ�T�h'���mX.�(8���o,����3߾at���Sl� ���X/3Fݏ�V����«����Ҁ�H���[��>��3c�.�/���0y`���?�s�t5���X�.���500d�1���[7[��V[7,t�Ǚ$8��y�gs�hŕbƶ-tiw��sve,C�^���!��7�����PX���)��9TƕE[AS�X������~	��3��;U�%@*f7�?�\(�����^gCۚ�$ ����d_Q0�'��>Q�ɯ��dC�����kD��?�vz��g��\��Ji�+:�z��x%�T��_ +�&�@9��2۰��r�#��_K�8�P��7��.�0m�w���_��/���'�e�Y�d{�䍜$gDQ{]n��m�
�s-@,gvt�\el�B��X�c�N�ݥ<͏����]��G��������L ��|�����$b�Tݝ�c�3��6~�dK�&�u�������ף�(Y_���o5_���7L���]�Y�1\��^�Ȟ�	ѩ,��?G:'��>��Ͻ?�d��M��(>o�F����YM���@"�'��T��]�e�Xμ<���R�� .m����X43.��im�!/�WGǙ9jr�|*O�|&�������O�(#��BP�����vp&"W
�6Z�#R�#��,v�-�'9K�q+3�C�wz��!�'�������o.���s��c~�:R�:-�3����Gz����4M��'53�m�&gJ��Cc?P !s�LL��M�4�Jsy�">����^��:�=��pѵl�)�:7?��,3�����b O��d�:��*�A	(�6�?xB"񤦟��=)^+��U��,�O��L�]<���D,����l�R�]�.7�����e��*Rp�<I�d`�s�d�I�8���|	s�xTz�Z~ .���I �:�e��C��%���	���N@�&��S� 边��N�r�@��n̡���*�F~�1X�9~X�� ��]�W���L���9��?nw:�����$m�q,��݋�r������,<��8�`���ш�z-���oy?Hm�\�<8�G�����ځ����3�+�{=�� N����n�N�� ��^5W#���5,�N4��| '�f� 
����3J�N�����E��.��%�⧰�q�E�߫��-���S�$bo�����G)�١),���Ӂ�M�bz�fe��?_+C�~ѐG^1FR��Y>w;rv1(�B`ڢ��j�ߙ݊6�e�g�{��~{�zTWQ�����*�G������kn�vLicU�?��	���r�zq�~a��4�8��CsX�w:��hR�z�8��u��*%����cg�a�Ȼˈ�D���b:`E�ϓ���*���<k):�g�cA�8I��n<\w��֤V<��Z?r��v�oy2�~wo2�W*�<�ꛩߘ>+��{z|�R �[��;��m��,�c�x��A�7�g�|�)�a�5b��6�p_��;������kPlOT��ln�I�nU<n����������`��ڊ>�ەG�i/�x뤒�/{��b�	�
4�q����
wE
��I�tȦw懟��Г[[0�nk�+^� �=bc��jP�g��wѬ�	���]�H����*6�C�>|;�����������c,��l��f�Оj�)���B5|>�����V������X	�)Po��5�Tb:؋G4~;A�������dc���0r�?��*t�"�ZÛ��c@�Br�vߛJ��{
 K�O��u.2����#ι�7tΘ5�A���$�?�������)�Iy�P#EAv�	����u�;"� ��}'��,*���z��<7�����T�Y��K6K��e�PE�� @��WbZ����� ����
ģv��پfXϰ�v�������ez�j`�B�~Em��{@4�Gc���)�I�u��ZP݇T۬2;vPOy���n�@pUzw@	��̼&��h����Dރ�wv��^�=)�*�w���� W{���h^-���Z'-E�|>�.CZ���瞧�/��她3�<�ł7Jk���5g ��,o�za������`��ʛ:�4������ b�q��/,���@��یi�@�k�$�: ��l��R��~P@�x�Ik�/{�ˡWd=��P�s�5����оy�߾�Kʱ*���}D�e�x�"���e�nO\�{<}m�zOm53q�MQ�i��.~��݄
�-�~�=����1:(���U1-��7J��8� �C�qO�� �0��oJk1(�g�(*߹��˾W��N����!.��a$�c��I�*�n5�BV��3#p���4���"&DT�@�c����q��66Z��>����P4�=��p���@�SF+ƨ��M�L�1��_�ts0�7ԐSEn�B8��?�A@"�wLm�V�ؔ.!��#`��:̝��������}���_��ڃ����.̑ˋ���ĤO�O�r��S��i{��x$Y������>o��ҽ��l���m��uL2�z8.Uc�D�<.L�9�caVg�( OA+�/~���F>�^{c1���3>���Ը��P`��ǫ	]�j6�Ԝ�w��5���ݫss��z0��8M��LT�K�ۿi�߱�r��# :���Ƅ�v���>5�J�R_!��6h�0���h���X��|$��b*	�M��f�/3���6���U<n�F��R���u,I4$t��n�
7Lyԙ�3�"m󤷮H���,��R��@m1�o/U^�,|j>��"8*�
M��hsaǤ�d���pۂ#��/��X�v�9/	v�V�kߣ۽8�h&YC������=��w�M�X������O)�[W�k�����,��s�N�Zw��!B��
/���v�J�e��ƈ�!��%�b�fmJ�j��xE
����7�M�J#�
y�8�c�\:��(�����T8��lM�8
 ���qv���@<�S���8 ��7��7�[�f(d5p������ϧ��o���a>��OAPcZ���`+�P�f/����? .w�ߘu��}�佖�祡h/��g�?}~���q���!�X\���iv�����M{���� �d���k{�����
���
��kl�Р�x ^�WK�#��0�`Q�RM[�@00��0+�$����<:D�d��vlˑ��� �T��@^y��@����i����@^�����Pn�3�.[pS� � س���W�hۏ4T�n�������gp�A:3���(�������d�{����S���ỹ� F�%;��-7w8y^(�yV�����h	� �ΑK����a<��Ǹ� i��&Ĩ�����kl��d��8���_.8P�jY�9�Ϳ���?	hh�����-pa^$@��x PD�aU�]��;�N[��]%���
�tpF̽�y=Bv��A�Ї��w�����v�;��B��u������V<�GZ^='�Y�B���D���6� ��fS��d�1��4���M4��]���g.��9������HE!(b�L ���ߴ#3R$Q��;[���_݋�E ���ƤV%y�k?0�� I[��l����3*b�pkҞ��h2p]N<��ɿ��Y�ҽ��r��j�p/�k�"��"ܲApĀ/ۨ�kSJ9���o�����)[:Y|7�P��B�6   ����?߶�򛰵���E�J%��qb��~B�/Q� #p�4qo��jİ�8�F�1XwOe���z8��w�̳��h^�^�S6y��C�2�
���&+P�Ȟ��K]�.�U�fT��"����0MlCޫS9aX%0df����`���6%�:X�B�lO]�ƅ9uo�">%��T�ȼK������Fm&���S��7��E5�/3��[��:��c�/�`���/��w��L)r.:%�V|�n�����z���������mt�^���L`�	*il�
q�n��Y��nĐ��xc3��J���n��b5
H��'ɛ �Oype���%�,Q�J�X��R������5��6�TÃX2��?�����R	�d3H/�^�S6*1�K|�}h�vԭ�R��c�7~�9���Ak\�n���>{���m�Y¾u��.mB����]LyL˨w\��?�[w��/����v/���`��"�d�ҥ�P�����e����q�?��0̠?�[��E�1�p��@��]��K�w���.t�f�&IoK����g"�+[V��5�����<t�y4�d�3�b�����uK[7~���k��g�2�����:������w�5� ��G����������������_c^3� ��J�y������_��E�ڛ���6��C��%�O|<�oז��r���,�?�aO���6֤�˒]�s�C���4�(�ZG/&���X�:�f���-
3-�R�I�W71���v5j7��਑Þ���C'.�B^m7yl��{�˵?�n���,�����9�ܽ[�s(�ȏ�<�Kcm�I���xfs�~����~Y��;���c����.�E[���(��6���y�3Pcs�#rq���d�0u^�B�����}�����7�T��p���W9��>�P�W#�R��af�o�,� vDxs�waQwi��o�ǎ�m^Ӿ4<�D�{�9�U�N�ouj�sɲ�VR9���ț�6����(K+�e8e��k�7��n�3��BԯJ�����87�x��D@�޳=AAqHG="��ȏ����uQ����D��d"}�^�cs��n��)�:� �%ϴ�:�T�4=�4t5�ƶ��|���|�g��w�nZ4H�s�^�2!��O�<ʑ0�ԭ8��-��iz���mw����^#�;�x��,/}��qm3�����j�!�_jD�߅Eg�SS��jc���jsH�ѹ�Q�X4��b[0��#�?D�&�of��KM]��G1;~���s�~Y�a���
�^>q��;��84v���z6��3��=���59=M�72���h=��j�9B��&~wM��U�K	���ٵ*�g�W��v����V����̬Y|��7�.�vQ�'˄���G֙EJ���?�L͐]��^@�+���;<7��a���E�2��w~"�c%����ˌV׺\P�((��'�r�Z��b�l�߇q���qo�oq%�#��=S��2��v3�J�A�!��*��"��q�k�ʬ��~#���<q6�@ڙ� w�ԁۖ�{h0{Ű���(Y���oRE���;[zyG�z�7�v�d������p�-�:m�҉иk�?U}׌�D@n4!���Tz]+
��H���M�d��u��J�E���p��i�_Z7�9(�9�S���l@���Y�ny&3,�-aZ9����[��p?�y�,v���g��(E�%�?��k�+������|W+!�|x �5�N��'����ŕb��Q��B�.U�]�2�������7�!6D���9W����lH��j��Z9�F*z�85#ńH�(��4��?��ѽV�zJ�k�
۷��*|KU:-�D��B��|��u�m�󙀳 u�,9�9Z0��U��M���R��%�&4� �	ŝ�|�<��*���:�ۼܑIs��p
r(�ĸ�몜�mb�W~f��>�/e���A55�$��¥v�x?Af^�j�Q:lKD�XR���V<ݿ��BP��tQf��a�J�����m���
5�ʖ6��I��BJ�Ⱦ���R�P	�P)ʞ}�[��k�dwqm�~���]���<O��<�{��|���y����o�6�6ba�.9���&����e���0�Z$��3��je;k6�Kl��X�?����55�ܥ�«'��Kf�r,W��N�i���ͷ&��k���L\�����7���ǲP��?y���4�0�D;���y�+�#�����ƫD�:�X����������Y4F�Q�J(��;�j�����M��-��:y��qb�a�H{߿�o$�+�KzM�-QtM��w��n�Ƥ�5��UD}ll�b.�Ո����kRZ��P,�2��L�sơM��U,��D{�� s-�h�;��Y�c�H�"���bQ��;�,��j7�5ʻ�]�w;�/k��wTM�L�s��zl
��t������] �K�S}��_T|��ܓؗ�1�dd���?�=��Mm��ء�T��5�(	�Y�@�i �;S�_ؚ�!CT���Ua��&���°��:���S�h�Yev��J�Vx_Ul��S�!�Ff�vOms���4�ԧ�Ш�9�a��xZ�X�H�s���f����1S�cv��&ʁ���	Ղ�>�Eɬ$b��U1��&w�R|���n�$ߪ����`߄�C�� l��&��V0p��2-f�|A�W3������+Y���J���Ҋ�.5��=<aLq:�v�Z�&u�~`n>�i���Ǆ�NF���XV@}�����j��)R��U�ַ�Z(�r�}�@Ǽ(_�x����)�\�}�6
K�/�:M��p���L[�H�C ��oQ�`N�V��\�᳀/AL���wiX�\��V�W����"L�S@KF[�\ �%"����/xQ�^�$ `~�����L��<M-�HqMUZa�������V��\�k����u}=DQ����~
B���i�A�9�����b��c^�	C��l�VӍ�t��rW�8�~�2���]��d�>k8���]�6#��YHu��t����^���:9c�F�^ڤ _�����hN�Q�uu�h�����¡�R;\�2mc3�F߆���4�yg��H������s��<�,P�����W��*G8�Ԅo�ų���"O*��e����eq��KDԈb~8w�kF1{��;/�X|q�әj
?�����`m�@@0���3�7��3�	�b�����_��������?3x�1����ѻQ@Z�(H&�Kз��M�n��1�����|�L�˃E�8������!'z5ج#~H�w���M)�u7�7C����[�'o�����uFSs_�`jX�d"
��P)񒶷��///@d�Vb
��	ӌV��`�xn\�^�C�<n���t�8�4�N��Y�:�W�Au��ڝ�]�R��)�jX��sFU5ܔ�W��Z@�IĹ�Cq�\o�����qV\�܆z(�9ځZ9��*�c�.G[����`��'��F59�A�Bt�����k����fYi�޹��o ��U~4#-�N䣘�R�͊Z�,�8�HG�P���B�,~�V�*A-�S��و�4Gr��o+�~��v>���%p:���[����~I�VB��y���Ft�F��A�L����#���l������zR&i��+�O�����@\6Х�xO�ʠ�"����pK�6/�0S�r�罺§w2Z��k�n��!N�u�x�W��(�W&�������6��P�t��f��<�����L�����z�<�8�JX�\�[��;���쮓t�s�U�4}L���o�pܿ1��Y���[�FF~�x��4�6.�l�������x����Jt�v�T�p'R�@\��g�@�x��f���z�F��y��A�1���;�j�%c���v~�����{�~�M�YOR��S��Z�	#\�"����rfh�}�hj�i`��oR��6�Eʸ�"1�ҹ[s96���$��OZ~Xx���I+�p��;��V��g �`WT+E�b����^���Fr&VH�*���|$��b�I�~JPw�#e��Rh�\OT\܁��B�11�j|��1s�rWtտ����>@��Hpz9�i���U>��e��dĽ 	NT�fƛN0a�ʵ�j���c�fO_(з:�$F0n�*o!:5!�g�t�%_�[�ZLe�ۥ�c�rϟA}���-�5��/�)��1ȟ�rkc��V?v
��+%�G���H���&��(d� H�F-���[ǜZ+��YX"T ��₳ ���D����!4��K~�LA�3lf��$&n�gd��k��,V`B�������LOv�1�uL/1q~g�V��yP֣�������G�� N�X�Q�c��@K1��+�A�-O�U8Pر����y0`:)~��d��N�>��fe��k���FQ#VyȂ��T�VP��ll]�!���u���#��x�Z�fy�)D����eȮ�a?6Y�r�.4���C�iὂX�R���?���("?�~���S�.G$��o��y���f�5����:3SZ'ԩ��פ�b��6h[�ܶ��3�f��At6��(u�k�� rg�.i��E�t%�ƍ꜑�T.��>�H��s`�)�En��tN��Fu�=4'��8��*��4���\�>��'�y,����F�����Te�y$G$6�=��H!̈́� �˜�൘����e/4���jZ.��˅p�����+T��bўˡPM���N���yw�����
Uq�q�wW��C����ܿ����#�Ν��@���h�񕩪\�D��
��eo\ܙ��Ƣ��

�6�b[Or������I9�6�@�@�����@�"�7Q�y6AVAf�ys�㞹.i>�;`�(�q�ڍRMd\ʀܨ�2�VV�Ke�����SK��{�S�����d		�ƙsx�鴇��-�ɼw
�*z]�}����Ź�a
��kp[��?�Pe2r���Y�
��f/�!�z1��S��PX�Aisb7����?j�z�Ĺ�@�,cCn��׹�������`���Mqǟ|"����f�����2�g��^�s�������b��/��M���8C�- �̯���Seݮ�?���?B�}�_��{��8���  �����6Y��ŭ�Q�5����\� lg��t^��L��$�)�|��:�fj@wVBWd`�g��U�hn��(�R���� .gR%��Q�O��d�~�����`?�ȥ��b��%�tDN�\�dOߞ����ƙ��ȓ�����������:����"%�ڢn��I�'�F�.w䴆_������\�����7�G�#C~��fr�J�:��u�m��{?<e��jG���~�vm[�zltA�X:��j�s�nW�Fr���mɴ#}�ewI�k>�a�ϻ�ϿGn������Ѓ�;��K�^c�I1�G��h
,%�k��\������( �le��\S��ڭ�'X�����&�2��%�FY�br7�|�;���L��v�p�&��#�'��Lk�O�Py����;z4bXd[��̞�����+9w���TJ��'�1���Rp9�:�6��[rw�?��G~�W�W��?Ż!FԀ��R�L�\��Izy*�ea`�)�t�kBN�^69�a��Q�n5m��skc�45�R�n8�ޣ�?�B�3�G	���$:Ɲ��e�Vm��'g�<'�^�>���ѷ���9E]ޢ"�[��ߠ|]	�-sɥ9��$�ǫ��4��3m�R�'F�'�:կ�4dw�|���[���P�)�T�CJ�]���#��[�k�C���9�����	Gth���:�s�Ĳ�����XWԃ<V{����ϣeiN�af�w�\D��������yH�� V钰>�C\��� �Y(�Ny�@�9�XE��3�x m@z���&�"��]�Y0�p�c89�\���Ε�O|�*^�Oy��x�a�l�	���i�S�{A� ��������3o�)#d}�\�r��#�Ȭm�W�vPf3�A�	��0\�G�������Ƈˡ����Y��S��n�_��[�d�jy`u�s��3SN4�y�Z`��R]a����|���xJD�{R�/���1/�*`�1�����lk���5�yxo%�tU�� �S������3��FHص���h� c'y��������ӌ=MPl�;i�5V8)�#|�"�떳���{h��;�v��bg���� t��,�K�B���ˌK�Z�R���܇%��Ʌ�:��M�U��&�!�"���ܐ���U���_.�--T���ڙ��,�������/|A�kתr���l���>�����̛�S|���©"&�(�:�xK��D��iHH���R��n��a�=]�����_>��j�����>,����U��|�{���x���O����t�:ک�\����	{���� ��>c-E�qc��}�������KߊƇ������IqI��V��V�s�2���߸�s��Fw���jIMߏ�s�Cj��������*�[K�[Ϗ\��+We����~�ii?�,^�s�БQ*����`y��i��|���k�v�C�iw��3�o����:7�Td��q���5��}L�.A%���<��\��������:�˻17�=��A�(���"APuߠ�����4@N��UQذf��f��S]6�y_S�a���"9J]��Sk��*\�Ȧ�WO3�awid�hR)���L����t���Ɖљ��<���������B�!19�L���ʬA'/�cx�{���j^{{�!a����
볖�)#����W�Nc_�R�W���a�A:b�̐oκ�k���A���[ŘR�`��s��l�֢��"�q��Xg,� "�-�,�&�e�2P̡�o���8�9K�e-������ľ>� dЌ��]z�5��ؐ��!�7��\ʫ
�0q�[^|ѻ@$��}+�ڧI�;'�A'�O)F<����_�~�T4_)E��M��>~���0l�L_��pu��9C~�����Gy���\����ƭ{X+ٔX�@���K��,��Wb;a9W�NhK����*���'�;b�2&��_R�.'ks2r�56�˫�;�5#��G~w�֡6�B2������x�
�ƒW�=�b7�ڽ�J[�5H���&���(5����>?�4Vh����{rO��d5I-K[��ܟֲM�7������YS�A�Aw�+
o�֚j�na���{|��}�6�0���&��d�d��q���CaQ�~��Q	Uf��4D���{vŠ o�1�'
i&�.cQ��n��t�o�ʉ�O���(���ɫ�63�4*/����~�f��%bS�J�Hj��{4��v�Q������T��C�Z����Vz��0��-��P{�֥�%����y�*���j����ZOk��~����jk�А�ֈj�(@���xv���H�"�ܙ �=��)"_1�,���q�ڼ[�|kA�\c��]�˃��_����;*�z06zȓ��<����WŶ� �Q��3q��$�r�M'Yo�VQk7�zSsF������\�'̗`����_M:RY������n|s��W1Nt]��4�K �)�i�*������'V�#x�b:P��������	M���P-;|�|�j���lF#�>��}�N��iY��%+�/bpsG���w��i���d^�v���Y��	Z*Nr��~<��D�^5|�e���P��'XN�[w�{�>g���jp�*�DG&*�N��!�����z��	T\vm����c׭ڼ��|�� �zR��0��I�`6�y·1�����3���Ip��7��`
���q����~���r�����X5�g��9k�ņ���o>]�Ҫ1�3��gY�n�"�19��6��F��*'�_�>oR��%�K?�yY\Ԭ̝i8Ծ�OcP���}�W��m#������|����T�����Y�R����wc|j���zF%�J��;NNUe	<��L_�$l-�a�iy.T�H��Խ�N��]z(!y,]�1�WeP��pV��>ڕT�١�HG�hܦ]
�nƒ`�	t�\/�,�)��l��W����%E�c)�E��h\S�k�a���̛��Z��Z�xd3�P�mq���Nr��Nc�A�c˱�,�VJW���9w��@ޤJ+�]j�Y~�R�㢟��C��9(�!I�_<å��p��3+ߣ�!���q�H*Z��jM	�h0g�%"*�(͉�$R�s�V��{#^��^N��G�r��~�\��3b?ΨKw���HmH~u��U���5�5�O.r�]������,E⨜��g�,�%�!�ʺ'�+�pn�×h�D�w,PںI��<���H|c�%[3J�|;�����\gnR	vJ����V�H
�6#þ��GoU����"\'���S��z"���q�<܋��T8���`�EzHQn6�:&��C�͖lǆ��O��ݪ�����y�l���W�-�޲�دrq����?Bf�0���S?��P��9�tD�8�}��%���q�s9j�dɃ�[�X�������P݄��.�D��EYM;��3��ѽ8���#�����Y�PJT{�x3�+v7JJ�����;��5���g�4����a~���%=@朗,u�w����1�MWŮ���ѕj	��
ot�>
eDޠ��>���-�����\i�}X�hWoIR����4�H��L㋏�Pa��3�r���7y�0�G������2���#%�����*�3��ɪ,�n�H>��[���1���El���������R��Xy��":n���oo�wN�\����[�?E�xO�ڛ�-�פ�W�D�MԟmQy�3pf�>/�l�A�x�g(�cz6}�2��t�CQ�� ��VE/��D$��dGN.��z3b��Y֒V�Y/�?�����Q�t'���Q2�\�
戤/�x�'�E����;��q��G���1.���9C�Zu܃,�W#��䯏wU�w�����mZ�
�be���O�i��{�&k�\�9hK��y�S�X�&����8)�<!�/h��x:���#V���nbuZd��|
N�E�8�u�N��ب@�xs��G5�Q��{/�b���r+"��;����8`�\�M���'����4E��hSo��o��{9>�-@�x�P̳��1�S�^2i��,'�[0e9O��cյ��ɾ�T�݁��(�-�����4p����5¬�nH�䙗F�e\�Ëw��Ji��������3�u�&[z.�VX|�m�;2�pN��&bH=�)�}�^������5Jj��2S�ac^��Ɩ>���?	g��C3�A{�5�)=�F�5Cب&��V������D�L9��k��4��=<Y��Ҵ�)G��)u x��ވ��>��.C�L��!�4b��7�Du+-� �������(�<^�h���wu��?e�v:��|����v��>S܅~�O�7����/ѕ|ƺ�;���L,w�z�M���D{��]Z�i.�J͡�������x�}E�Bk4;G��ڏ�ʁ_@��'�4sRyNM�u/�2hAـ�[���e�Zλ���}l�e0W�nc�WY�@ [�9)7\ɜ���ʊ��K�ca0C�E3$8)g�Kb�K�$�h=]n�=(�<�1~$�u���}5����u�ʽ�BAW�t�8[*�k��I�ً�Y�����R��rƸqo�s��ƌ�.l��KP��KާB�����^UCN�E�)�rhE�u~������TM;�`Ne$��>*2 ��k.E�E�8Xd>�7��ZaS_�M�ٿw"�B)M���k?HL�yW ��*�5��D�L�|l&���N"Pj.M5���2�X;���y��M��Y���Hޑ���c���j!�Ŋ6	�2;Fms����RA���<$�/>���r��ċ��H�r��dXT#���+2�9&�+~�c�0RJu+(sX������a���J������O^��n�W9�l���ف��w�_�tA��Tn��_�m�x������#���>��[���y�i�v�Gh�+u[�>V"r���4(���q5IMVYs�%b��`Y��r�;vX>���V��dx��`K<��k쟟S�s�Wþ�3� �Hf@O��Vw��U�-:����)�=���c@?��Ar����n���f�pN���]	��M�cfr'ܮ_3�5-�U;�;��G�2n�Ug^��䶴�/	KX6D4��_p2�s�C���H�J1�����y+��I��~�H�ے_Uu��*D }柿	�C�w�� c�̜A϶b:4("a�{haU��B�C��ϵە�h��:+���;��@FB�����G���]�a�(�����vҼ׊F������?�Y����ӥ;��ɍtNZIN	���#S�C�V)�B�O|6֏���E��U}�'�rx��ǞO�Q�;��u`]�zvu�E�p-��������;V�׊nbM}@S9j�,#��V��Y��:vGMџK#}3��b쐨D��b�u� �ʣ�!�l��w(v
^��QH�����=yKV�� \�I���Q�� 	,��I�7SX�Kg��n��Qуd�����R.=�V&�u�:	9}+����!_6\Q�cݘ�O�Z�����b#��b}�\n��t��L�帋>5�ƴ��p!�5��*��䰺#�T��`�2�<�b����1�s�-|v2�6ND?g
/6��"�h+O���e��˒��ZQ���-3?�9j�ʑa����1���G[�`�m%M����X��=�s�nNy�����v[��z[��*��T�����lE�T~��;�KP��%r~}��%t
 䃆��!n`���Vڤ��r�י���; ����ٲ����-N�F�\s�I� !D���;�'�0���W��$�6�vG���
��I��P������+�o&����N~؉Uў�?
'�,&��V
!xՔ�'\�dU���X���XƱ��� d�6֠�X*�E;1�R�[R��ȹ�g��f�![���]�D�����εl¿�1�x�X|NQ���꟧��-M�!>L�?�|?2\��G���L��k�f����;~ћ�K�I������^e-$nWv��m�鶵q_�P�����'e�<�I�.;eǎ�-{C�܋H-����e[�-�Y?�	��v��su�����ׯ����Mc//�䱗32�D�>]��á1�h����H����G�b��5X�3,Y�=X�/����Q�Kf�0ӭ��e����W"��z�ܟ���Ũ�I��p�����1�t&j)��^��E�(^����ެ=w�G�=�i*��R��-��E��}���G)-G��l�B���<6�x�����~U8��C�pv����S�K����`������--1�.�K��1�gPfa�V�����53= 7H����)vO�sd��I]l�k���k5�s�%�w�t9�B���Y�[��l1����ɞk��ac��^n�A����7h�blV�/���b�V�?��>2\8�]��Q	Z�s�Myj�ި���b�D�5�Ǘ�����n1����$9/�q-��w^z���Arx�����ݳ��Z��	Q���R�q�z�"Ӹ���h�HwU�E�?=Ό�;{����K��:Wáq��F�L~ɒڥJm#�����s��|����࿨r�ԝ�e���
1��z�uQ��{n
m��,{�fyF�d�r���1�0?�����]��EX0O]��{K�x�ci_)�⺱���k�,f7d$Jԭ�����g�J�D��&K��nرn��8G�Q�M�u�>�2� ��S�e��ײ��X��]�:�?,F���N�/H�xL,i�١��i��ҽ��L�53��]�бīt��T֐�����̏~U�Ut�������=��}�{g�p"M�t1�D1��W]_�?Q��O�/�R���L�nmٕt�p�*�Rf�JT,���� !��e�0����e����cӺ^m�3+���?me�*��+N���? �e�1S]#c���ެ]���d�K���Xb�Y�^�oWr�x��쾞zeކ�����`��R�j�����e��J��i"�T�v+���%�-K��OmȬ���q��䑒�-J�����ǘ#y��ړ�9(���a�Up��.G�L�.��h7X<C&���11z�މ�߇e��?\�^|�l�Ē�,�%.���G�\�X>�l���1�ǃ�ڄ�>C�G�6�z|��hG��<���_��U���e���B��dk�B)���YY;����VpEO�:ñk+�[����FO��'D�<�wk�"��]�ٟ�1@L߇n�̜��qv�p�55�@�Gߓ�	aPKC]̊�3l�Y~�o�3^o��T�ڔ~I�T~lm��T����xM]Y�d3��w���n��.l���/���8vo�o��)�~q���"
O�6�=�h��|������Q��ީ-�i��p���zv������F���npa�Д��%����w�����-G8��BT�1rz)�@6^����՜T, h�u�*R.��ͯ����A�i�n� ���.}���6��;�dY��4d%Ir��7����t�/�]f�����z���-��?�|��z�2y.��wh�]ea�"]䬭�����$�I���c��ĳ��ʭ���u�7U����1f��W�V�x�DA�Vo�,ߝf����O��7c�뼄��o<�=O�;�\��K�>I���A#!a9��SC֮��ȇ�����tؼ��EP��
��nj�+;R����H^ogo|�4�A��x�ɬ��R�&_Z�쫳��������H�}a�ʚR��"�t�ȇ~ZG]E�ԟ	K�����s�ȑ��"�Y*�[\�UHF�"X���j���A�R�,X��3�q���*ƒ�p���U*E�y^�$੩�A;�s�;Ѯ~h�y7j��� S3!6s�
��M}�c��Qʺ/݌|p"���fT+����9<&@��*�Ƣi�l��`�w7Z�(�C�{Gl^����H�%��c�>{�׎)'��!Ə��N:%�s�;W��63}|f 8y$�F��X�%i��m�j�xo��+MG]N;N�eo���Q�����!x������ʦoK��ܡ =%��a���;:��ۿut�������'��q{��;����*(�:t�W俘��q>�??g��h�=?�&c�P�$�w�,�Y�S�Te�zr�*ƥEa�8��}*���u`�m�I=�g�n=�1��p�OW������k3���O�#f`.R��h���n��紼�L��>M��|Zs�nތ�%�����57��c4�R^ 3��9
���37��oEmL�!�^�(�tQ���!�E�#
$���]w���N��V/z���,~-��j�� ���ͣ� g�͔̈qD�nQ����á�Mj���j@�.{�EL@mм!�1EY�MS&"G5�����85���tՋ�¨I�	
�پ/�o����9YǴ�r��5�{U��>�H����1v�-('���o�aKs�`��`�E��r���m���t���[��ln��)��nW�#c�Ò�Egѵp{�ô��ؒ�-��zܢ��'@O+�Ǐ�����TmEAe���n�L����w�>��s�����G�\!t������>�!��ѓAU"���[f�*�Kq4���1M���,J(o#���E���eǦ�)�8O+g�G�OSs��Oj�,iG��x��ސ���૟֓de�OY��>dc�2�bÕn�U�tȊ�Y?����8!��>M2�_����K^�{����I����Ȥ�FW9Էױ!C4ҷ�,u84��u)���}�[
6a���{��vq�����)əmb��}��r�ec�HQÖ����&�ǅ�|�4X�:]�"��p����i�<��U���lA4��p�Jb���2IE�
wT}�N�(NcmgP�Y���o�(0��0�Ø�|岥�=�=�|��=2�xf���{:�����C݉�g��RM����yG㝨ޅ��ɼ,�~8��	����9A���"��ݼ�@L�!���˝�}�}̑���hɼ�	�`g/Q�+�0�N�<��Q��m���{�|4j�
���l<ґ�!�yd�>�_xR�۞����,�,Ag������&HB6��V����IGbo��gz�l��� UXp�V 丹��cp`4�E�͋�
>����`��5���6���<��>@�@�L��
��[/$�l�Ó$�5l����䵠�[�,�3� 뙷n񖎋����C^�4u5ZR6*�����?�B�@ �.���_����H����N��w羨�bb����K���O.^8�����p#F�]�J���""�P��꬗�Q��Bv|��1(j�R�dM����!�\����&��|�H1I��X�ՆЙQ���K�
m�L��`��Q��V*��0���K0��Dex�XCM4E��r���J2��n�{��K����1[Ϳ��哆��M���b،f#�6"9��.�Ab3�K[b�d>�?uG�=6��:����Э��v�U����NI˶� O�ݱr>�O�f8y[�ЀL���c��T5�g�W�Xo���[p'� ���&��r|8e��,�߱�� J���Z�j\Q<@d�8����ӷ��"�߰����h��j���Jl��˘��}V��S��8�`vRu�L"f��_� %d�%Ǘ�+�[��r�����?;:��4GE�:'��_����O3��ġ�	�\`��[a�ۖ�R��� ����u���&�0ҁadpI�WZ��VڣfM��d �䥰����I	��mx�1/�����G=�"jp��`� ���Qu��U�W��)f�����а��ݻ��5W�A����ڪ(��C��+���4|b���TϞ@'��$�`X]
��--ݝhg�v�����VS�IW�Z�w���V�:�ڋ��}
b��	a�Ӿ��.\�I�q�t�`?l 7|�&n{��U~QF��*���&[�,r������=��]Wj ksw��`�y�a��3�9�b;Yf;� ���O�	���1��W{F) �g2m�� Lm`m(�ci�=z����Uzz��<��?��䄚�Q�s�B��,���n馘�{./��[l���u�є���d/�KN+�46��jW�*6�rM�^���x�5z�bG|{�����`ׇ9aǜ�G]��Ū�Y}�.��6#�VSo�� �#��M��r�I;}A=�Q��0v����I([�����A�k�hVD���]��1{k���M�:}����lR�y���AA�u��=�H�����,(b�̺ӊ�r͞6G�(����A]�o7�n�b̺�e_�5�7�I���;��#��!�-Q�ަ������(�{�6C~��m���XdS�\*�	ˏ�(L���_Rs�\@}��`X7e�/��Z�p�yшF	T�HП�d0!Wk��q��P���! ��M�����	Eb�57E�����f�[X1j������&�PY�{ڰT��Su�䞇N�c0��6��>��l�f���L��a��@����N�#{�v��[!8���*�;�DΕ4�hU�E|�C�T2ѻ4V7�=��°�Ǝ�)S�d��G�GЄ�Xs
\mƭz�%I���g7�~9�܉O���-	`>����h�	��:+1Ú�@R��I Q~��?�~Is��e���;�ݥU\��9��F�A���E^�.�W�$�[�¿��2r~�J�;�?�:!��	A������&G�Qx�EIZ.)���`/&خa��YE�r���&���eW�7 .�� p�� �@�t2�n�fy��+e�«;
u7��$aW��p���BMzo�K]����g��T"�P(v~�z0Mw'��l��o�!�X�;~"\;�N=)�+)�#�s���2��<�*!����Y��f����T�!04�{J�`,i�����B'��uL�@���~f�L!��&Ͷ{x]����-Zs`���l+�
9X^��5�\��$���?�Qo/
�] �q%WuM����~eG�^�f��U�T��qƑ2%w�ى�J��tw.�ůK�]�#E�-�c3/�E���9U��̫�L������|��"P���B����ECڜ�#�N**�l�T{M�D �"�U��j��m�$::���~�NA��ċƨ��g_^�|�\��Rۿ��9��#�2Z	!��^M/Q�Q#��dz��n��f��� �%�)Pv�F�Xj��d�O�b;c+��0�ՠ��ler�ho��*����#S/`����C<KG��Xg�`�#��ЮW^Z~��=��6Z��{���Ŷ��2W`ji�ԵLWյ���(.��ۘ���h�`^�׎�~��7߉��\�"&Ѕ��׀���x5���WM�ךLAޡO�[�[E�/[�cjV�.Bf�6Zp5-T�̔�""���w��8�Z�E��a|�*t���v%�|�v��I��z�
�،�'�*�EO#�<��78���{�Vr��7t@�F�\`�Z�_TE0@�i��w��/�
��B���2&|a��ŧ����W(�NY6;µ�R�a�8��('�#a��ՂH���� rd�$�2�m`�E!��r�%�6�})�|_��;�
��'�[�#�!d�~��R��\C8ƺ*�~��`߹~��6��W�
r��&�;�Ծ�\w����/�g|����K�ĳ���~��t�ɉV���/��=����@q����v�������i3�w[�o��-M����5-h_����3:���p̴����i��ϥv�XT'� �h?��x���W���p�k7Z�I��4lc!�X��x3%�-��Q�Հ`�F���������@��_����l��By�]i�a�=iF���,�h[�*�D|#,��y����̍?���dV�ykߍ�	6��b8���A�?7Zl��$C�������>8]�g`��}4~�}V�R�K@{�k�TT�?77Є �6�fʲl�.�@mxSr�Q�xIL�Ƅ��M'�/}�r����X��r��iR'C�6R�sP;�aÇ�>� �0�{��P;� X���&8�E �F�n2�蒱��:L��@��u��Ƭ�:��������v�?������F�`�N��)�f�<N�)[5(��ϟQ�~	�"�f�(�V�-�!�۲�c�+Ńl�M
n��➻�taq�P	Ƿ�@C%�moڠ�t��U
R޵�.��{�t��&V��;�G=���n��Kͣ,i�k�YIM�'s���R�{A�V�k�H�T��~r���&T��"���%0̴ ϥ�zݫ���x&b�碦v��~�Y$Q}4�v@�q��ǃ�-o�����<�P]��ź�`'k]���A�!��D+�]x[������;<����OM�'�3c��ı����Cs��h����ǟܹ7XȓrX2	��,���%� .*�q8����� :uO����0R,�;�����LN�6�OpĶ����>��2��˝�tKf�:Bg��{��J�T?͉�Q������S������0���C4�
�Cc�7�y	��#�{Ba����/��x��+���k�Fy/i�`����y�DE�A�1+�mBG�������+�|��H�R��-w��.�u��?���B�YD�/�S��ʜ��L�{^����3T�?�/�.GI4wd���ೲ2HB���4�/�ލ�����%Y��Gɀ��2x��7T�Zi�s�p(�A*M��0
�n1<5"�㴥q�� ��)1��]>{��$ġ��5���o ��<d�?ZD�z�aDz�i=�6���?R���4�Z7�`R�z�z��:-"����}p�3
�������i%xe�E8�A��/6Σ�-�_�������ǟ!˟ݩ:�l��Ʒ�]�N�ѭ��\[UN-���
H�W���_��֟Ӱ��K�`��0n;��k	��oCT���X&��[=.�<��������$�zal둂-�^�
3�2�mē����O��a�v�T�ኘ���v�?^���o%`j{��Q;�r~!X����MҚ�!^��x_��A��m�?��~���-�p�3����N��)���C5�I����-����a2m���_J_�v�m��p_����K^����͟;���Rλ��T��ol�uc���S�ߔl/��V���'%�cMsCu5�.Q�3�W��$Q�8S������մ}��T����߆Ҍ����y9������=�7=�n�*>�lC��6�۸�6;��;���-��޷�bY6���Uߖ���H����0�'4��#�W4�R��r�f'�_6x�����t͍4���E�zd&�zتɼ�WB�G��}C���Ux{��K���9��V�#i	�3�
�=�YV����َ�$�{�3�-���
g�kG�o���Ic���	��&�8�g�����xF��R�2d�˦���XW>v�?S����TZb ʟ5��q?��m&x)Ӎ��9�Yκ�E��Mv��7�+�� GP�܎x����ʫ�cw�.�2��&�7��+�g�<�h'm�w�8Qb�S�ė�g��(��p4���zd�a����=O�f�C��L̙f:/$U6���������D��_��O�zw���
��H�9�>�'.��Ĩ�A]�y؍ʕ�|��ɒ�Z[��(|{������ξ�����#�ʡ~��[�g��K�ۚT�t;�eKY)f��yN�}�c�B�?��2��K0o~D�y���Ҏ��-�z&kx�"�2�o(�n�$��ܻy��=Lz��w�??Q�U�~�j��[�E������-���f]x)�}Ӗ����@������'"2�û�4�3�����XbO���[ҭ�\HԽ.Xm�}��07���T�~��k>\0�����?[ұ��<���*9f��L�ts6O��<W���~~�e5�M�L�0'�'��ue_�m±'���{�+�FZm��\]i $�6e��x��sgG��58���g>�� �^��w��>�
F�����b�0]��:�:�:�O��ι���Bp��֙���@e��f��Χj+ l��g��,�	�q��)<Q�#}Z4 b�K�2���nb�r�gs<[���������3Y'�-�*�pG3W���=�7���`C7wu���\X�YR��e��$��p器ù�&):�8�iQ�&������z1���k�	�ҕO��t?��� �[Q���m��������=���E���:z;jEe8����[/�G2��,D���7=��q�rp����l k���U��d(p<V�������ժb��X�C�\�i��B�KiGfs�C��@<^��bϒ��7|(bS�zq��UE��k��@�8�Ù1g��<� �ZyU_�V�V����P��b�zp�����h·���n[�M���)����$�qbh�r�y���DW�G�N��u��N:|����4TK3AP�dxV�GQ
v8C_9~���a�L+��N@%)�%<}��%�ֆ�5�yBz�wo�[y�IEa��4c0]����v{!��ldĸG�7"�lL��i�Е�����8�ȉ��6�m�� ��J8�>��')n�%�����r�c�:b��<�^�}�R�#]�ie�I��HGIԽ�� ��+��	w<�,|L#�[=��������K�S�L�S��qEd��7��ᛧ	���gx����1�Q`�u&�Vփ�I?GͿ�2�}��7:	�"A����h��BH���A_�<g�ee���>������;�(К	b���1�p���XKn[�F�S�{���_�?z���8V���H�zQB�;�� }hf��{x�t�鵛C�{:[;��@��Ղ�)=�G�#
e�'�{ծn�=�;�d����pt�'��>���l�8�4�p0Eܜ�b�c�����g�/����eY�g�����wW}�Y��]��;A���C� ��˧.�.wJt銔u�T��2��B`�����؟���k{�ڢ�ޥَ������eVb�w�����)�/�O�5��?�z�"�W������{	��=���?�x�1��(��TZJ�V7�v���M�O������K�i�rs�9�m�>	�̟�����&���S:	)�e�I
��iяmeO�Μ�><�'u��ڊ�=�Y������r�F� ^�*������>P[b��2�
�<F�'R*��C��s~t؊Z�&'������Vҥb~� ����9s�#x'�_����\�-��@\�W�k��9�D��j@G��VkĐЋ��~�Y��v�����6-��8o�����Ȟ8��	m�Ԗ��_�0"-O7/�}��6�g�"�4b/]�0>q.�RT��D��ƿa/J<�vQm��%�<�g B���������GB��ľ�ס�]q��������g��eM]�v���~:r��{Yw��4/I6�^�z�g~!�W��[�w��`��>����r�Y�z������>��p��1�'M��eyʊƶ�A2���R_����_	��P|�S��љ�C"��R�B��$�3���\��ů3�.N�=|�T+FAd�B�6Xj<c�����5����{g��D���@�K�mpeM�g��W�< _�+�JT�u����/���lbn�m����}���n����g�m�����w����)���i���"��B'�Nԫ����WY|P�'�i��'t���w�sp�bh*�,�2h&��n�$4��=�ljm��( "es����^�]ׇx٨9� �/: �q�#�?I��f9]���ȎK�%��",�A�d�5qH���/�E"�E3`�]�)k:k
��l<q�ϫ����.�,,M�{��6B��#�yl���>�M�>�*�HG��ͷ�͑v�d
�/4���ׅ}C©O)��R���/h��/��^P�Y����f�W��F`�$�z1�:b�ˤ�s�ٿ���VÒ�9��b��k���_;���ہ*�
���*\*q��uRz$ބ��:�6_�}W�f���f�g��:�g��I7��{	E�Űj�ֹ��g"2����!ߜ�Q����k����S���	{�菸�����~�|�<�u���r1Č������Q|�7?������Ū]���m��3bg����-���9�lBBa�������=�ePq&A�߆1@�FPG�[�G��&|9�J?�&(2�h;�/�����޵�hO�f(���������G�&i����A�>�OD�+QVd\+�q�T�L�%{fo��yCƥ2B�#��<�9���_�y�����~���sι[{�i�7l�R���m6V���Ϝ������ąH=磨����T�c8G�A�X��LcsS��Sr��1��{���Dt�A,��u]k�ZW���;a�ᔃ߫��˘ā�T�?0K��$�������ˊWeL!�@b�u����T|���хI����1��ar탯{J�B��+����H����Y͙t���h�U	�oŨV�*�0��YM
����S˥Bw`��~�-4PUq]z�@)�7s�S`�p!�,c�Ѩ�c=�+�y��P��Wa���i�@lxj>��)ej�}x�7hQ�lNP��qQ��R��y�%�Tp��Nvs�m���bV@�i�<U�L�][O�'J�RM�����),��5ǅA9��*���ٚ�>U^5�����O�I,�5A�����1�#F�����n���:�@�t�tIfF����31;�9�0M�_�:,Z��v�n��_ �wHXn��	Y�%�0e4�-gݖ��4�A�ᾆ�ؤ�M�9��dr�w�����}��-򺹽�s���{`���V�7ּ:�l~J%:�C�4��bkdf���ݜ.���s�u6LH
��`���[�J�/�<J��Q�ĝt���ts�{��t'$�tF�ӛ'/ɢ�v����~")�:���� ��j�)@YʵoC-������~]硍�!���~k�	-��\��yBi�� �i��N�k�d�@�d�����Zݑ�0�4�Hb�zOt�͕GY(c�e�SML�I����K[���{m|�ۀ(n+F�`�Ԅ��H=�*���b��3�
ܧ{����֧WA���e.�I�ra��p_��i�s=���"Ƙ��&�N���`� ��.���n\��ӹp�kQ���e3R��~�8�df���mo�Yi��YC���垐#e,/o~s`�� ��+f]������	�h�?����!��\S�����<�y�^�=�n�ӑUo4k��D�)���S܎�Ro��oH/�7��~�������[��W��u`�R��~f���k40�ţ&���I��j/���ANB�٘��R�e�~	m5��^���:���r��0xx�^�-DS��	�ۥ�%i]�y����9������Gz|��RX�&������i'Q�׾�Y]g�V9�H\�6ZB:�^���֛J������t��ц3��ym��/���,0���fG�����J[�j�����1��Fg�l�=���)U-dQ3�A� ^K�#�� =�mU4_Q���Q*Q}o�kc�,Q,���R�}y&T���|�Y��G?)�n�j���%c�mW�}�����Y�?�'����L前Oe�G�"6�a����H{|���^]z�I���XK�v��9�f�t�Y�o ]��_D��������\����9�F�U0!�`2���V��_�������.3��Ҡ��C���G�^����ځ������F��+)��Y�<0 �,�5�W#x�з1
R�i3��/��W-N@NB���(m"ngH��rn5����tτN�.vƶ����s^0�7�W�d�Z���x��I�[�@�"�1�qm#�d-b�az~��=I&$6����1�{�'�s�dx|����T7|!~���T���{��}�dK�J���c�� q"������cd�[�!]57jt蓠�n(X]�ˉ��ل��t�������U$7YH����*(~(�Y�,���a�8�>��މB\X|�:F���K��zbQ���_s%5� �ԁ�|�2��Z�#e�O�j�D3�9'�j�[�|`�Vy�]����ϔ_��5�"�IVob��`'��&b�|�eE�^Ԯ�瘝D㼄n�s�/|L������z������� ��a��
�4KIa��3�0��q���9���m�:�6��~��K	}��ʒ���{#X	+;��R�@h�ϓɂ�{���o��2˗s<��t��_023��O�৞�9���(�ҜSP	 �G)Vq��	HE�ޔ �����{��6�Y������{�d��y��g�缌�򯙭 ��5K.�#L�.
Wd��D��XZçf�]���̕��Bpy]%�YQ�"Kg��b.���L�u�nΎ-]!SU](��!5�i�\��+�/��Z��FN�ʌ�`��n©�|�3'V@��y��m�G����밆螀�f�����Ƣ��5 %K����)U`ԋ��2QԢ��PTk��Fa-����f�I�=���#P5�O�"�ܘ�?��Z��j����Dtn�d�!gv�$����� �F�AC���.-��6o- sM�*���\ݚ�X�l�c�����)+�f�F���)b"����>�e����K���v��H"`kC�����57~���&�r�B�Y-H��0�Oί��l(º�?:I�$��V�[D�iL��]�zK_��m~`�T9�%VW�/|�XNx0,%�Jb����^��Wd	ء��f��m;����?�"��|ZU��R���'����\>bk�uQ ���)+R�"�:��]���?�@���.
�]�L�$�X���[/�����FK'�pn�����I4\�N�k��9W.��K����`�j�2N�̩��-�Rւl����N�I-为�ǁ����̸����V� L�ꀔJ^t58�D,;�9HY}b�R��9�=[c������N�so�ZC�&��-@w��,QC$f4a�;��&A�m%!��nW�L�m�Y��~�<3}`k$����L��S�}��|gS6�����K�R@Z�D]<<�\H�y׮]v0_�m�U�P� `R�BƄQ���?��'1jm���#2n�@����@�_��<�=����!�����"�/�u�$&x����SV�,J�=��
*j�;mF����BL$«�;�J"v�n���S�����1�h�1��r{��0��AII��-�,���Yz=/��W�-�,��;,�f�*�Ԧp����[�c\��Ȝ ٩b�T"� N��8��p����!�s���~iC"����f���&%��m����R�O�_�5~��_,%o~3��Et��6s&�mY
�L�#bn��ρ�O+]��Z�8�)���};��6���f�)��H���/x#��;9:8Ǟ2���E�I�����ր��?��%�E�?�[��>P{��/��W�R��,��'�F���zg�����5��~��$E�#;��9��΋��Mw@x'v�������ѳ�u�R�~s훫hG��U�ag7�x�c	�:b�]�i�_��}'2�\���P�`��O������.]E�XW��wߡ����HE`�!�ѱXvw{��~���k��w@
�,U� ����_��$f�ӆ_&&���ݠ�A/���M�����"�rY���[�R�	�6z0�{b��,��"I�Q�"�7�ՈҘ�_	Ŧ�/E@����O��5 '�����U
��c��k�Șk�����$��W@H�m!��qN8��ߐ�km_N�r�(� ���5�C4|ڔT9X�h�5o��{�C����ah�p�F�F�L�?w�����	����ŵ�C��d:��	,܆��+_�nm��깱EsWen�a#2{�o�.#sb��%V;Y��B�:?)p���{݆?T�/~�:ǋ9��;^3q߶2j�ۤ��G��XA=��y2�p�E$3���ύk��|W?�����gYP��;� �%P���G힢�6�_���+�&K�%�����5l�Q����{�E+/���9l���.�\��̂a��1<�6;פ������PN���+'�YPW�Ɵ��Qd]�=��W�A��^K���"2`uI �J�A>�p�JW�%����c��̍�W�#�nJ:ǶY@�l���>���*Zl���� k�w��2�n�/p^�x�Ri{�5}��0xx�F�`�N�
��c�����5"�F�ɐ���P��^�>�-����Iλ
H=Ǌ�7D�� n��:��ZlP3I:18���m�V�ѱ�X�I�o��W�	{�1x��nO�4ex�_�Z�����2D�@� /��h�2er~�@[ 2���e�J&���B tc��	+���uz�P�-]6��;tx�ى�SGP���k��Wt�sｺ��>�ނ�g�{8Pk��+5�y�jS�̋e�v�tb@�W<��Nh�<4]�L��
7H�+Y�AN ��,�i��+�t�4�1�Uv(���u��Oy��{��LXk�4L����d�>�%��*��P�z�b`��1_������u�_�y��������K$�����n��A%��<��r��tJ��L}�OH	�~1>`�>�	�+2Y�131zs�\bzN@��cL?�a�b������3�*WU7�8�*�o's�A5V3�>�s���q��?����M'�V���a�|m�gP4��K�~h�a2���>`?^@��
�B��tG��?�"�d�v�_l�;9�MO���N�ى�)������Ȱ9 {x������,zk|(��u�b��/�7��4d6�aܻZ(����<~lML8'!�C��y���nY��$�B�Ha�V�����^j��`n��&�3�s�}ß<��g��<��ˈ�	j�X�*}�"�
��@"��a��f���Q�/-�uqX���z��D`����kxACI,�����F8q(z̝x,�2(T$J�i=h6
ڜ�kuZ�ֆ)�85_7닢�֨����94��L4���
kQ��
����(Ӳ'/;ޛR6����E ��	S�:���;U��uA6^{$qn3Lt�� G��8���g��+�k+����W�w������܃�� �Y�IHQ/7�G�7�؏8�	YU�@�ߕ؋d9�g}�5�:3*ք;R[�D�u���꿜."]�����KA'����ϨX���ª52���%��Y3����4h<B�' hڸ'�3-]&�lA�u��X����z��<���%�TU�W��:n:�H����ǔ׬υ.*����'}��9H=��#�qĘ�#233�y��[���������o���5�x���
�nBc�n3��I�����׊�h���hS�c�W��-�a ����'W~ͦ1n8�%3}��S
�G�t�K}%>�^`3�B����&-��X�%� |���c�G,G���h�~�<R�Q��M�\Q��K^?o�K~*���N�Y�Փ�����2�9�?�3`��c�iG��_|q���e�A7�7����5��t������k�>߿�}+���G�=cd�qf�ɕ�~~�r0���b�	������t��#OZ��X8��{۵;{�sZ����yET\t~����*�ZX=.�~B�KiW��Dg\��/�� *$���I�1�aT�(�Eo��G�3�X���F��ײEU�3�o�um�o���X1Z�~}<x�F����7��c�5З;L��^���0گ��E�~����C�z�E�{*����[K5�uE	
�co88��'�p�rq��KF+SY����?I��w�~1�V 8�v	���åaF�E�7Kf���]���{(ģx�ڎ�����x&пbG����XY뢢J�S�4i���ג�tǱT�Vj�h�^��BU��L�~@�Z�or|�y��@�z IAܒ�x���>��y!K��1�clF��am$O�ۮ�u�.Q!�U�l���F��R��kh��� !�t���r!���4�
���^$P�ds��P�u;�9��_�pA��>)���~b_��C�@o�O��P�[�Eo�VhK���<�5������_��G���nɤ��{��̡Rz�u��f0�8�RD�S 5{�:53{&���m�2�F�{���,��i��-t*v.ǯ�
E�Tu�Uk��(�4��a�I�R���~�P��|��=z��_��FV�5P`$��+4~���1��k/���u(�@�Ϊ�Hv����Q��Vl�A�l�}��K� ����@��|�y��]\Ƒ����B2��+M0!H%��+��\����\��tX�K�t������?5BVyX�f|��$��(s�2e���o�����C8E����ⷌ�L}`'1g ����ԁ�Y-��i���BK�r0�;FX]���_�Z"�ɗ��X�Uc�)7-`�K�����ֳ�߲7����q�P9�N�4�b�2�k���ױ��������Q�y���A�����Ѹ���Xjd@�R�C�q��jݢ`T$��fe�s�G��4u�o��(����´<��aW+��"@�p�`)����f�	c d5�r]Έ���o�:�R�`�x�U_:擾t�?�RG���%h7X�E�Y���<A��V�;Y��KVZ֧x��3u�+���:�lIQ��3�|�G��
�=��&J��Ӯ-x:��^wx��݂���C�C��)��Kt5V����Ez��n�*ǯ���"��M�M�W���<be����-�i���qK�V��y�2O«���u���6�r*��Ҽ�\����ڱ+�nG�c���.9O�B���y��!�Н��k��q|�
�`�:�	uW�2����6Vt+��~f���p]0Z�%�M�ۑ{.ʌb�%�?֧��
2{�,�+ �~7��Vl_$v�֘;���ҙm-��7�ƈя|�K�}!�^˫�B��@׆0�b[x��t�[`��4FOx��/� �}��=�B�5C,o1�{�rӵ�3#~#�1�?���Q7��AĮ�X$�T�m��Z�`"A����e�S�f����2H�L�ÝS��H��G�N��	�c�e[���Zs����O)�L����#CW��[�v���b�T[u@����, @����RŘs4�/������Z�z�	Z�d�yk_?-l���z��&�o��U��f��Y��	̡��T�*/��G�f���+�0�/3�y���:����AxX�?U�X�9�N�	$�֤��h \�2U�Z�I�eA��+B�TG[�"i�* I�����H���.j�Q��H���]\Jz01����}���N$&����z�]4j����w�W?�! ���W�+��N�,����\������RD�&])��/D�F�����j�a�ZO���枈2�E�asMt+?� k���ji����T�x8��@kK��S�?G�a8��7c��Lc�����\��Ȕ�
,h��@uF9�e+�+'�d舖�u����V��nS�D��[t[�5MIԭ�z��Y@WZ�$a���I�0��:���{n7�,��5* y:�"]����8�oRPpw���`w*{๡���e:Ѥ=��������Qy�&f	��Z1�E�H��?]BS�:2�� �"��t�+M���0^���p̥�Ųb&���0�M��'��܃̅V�Tt6��0B_��ΐ᳉J�����T�Q�b�
Ѿ?��6M!0���2��tb��(�nE�c?�m����֔D`�[��^�l�z���攴d�0�c��!jf���ǽ�32�WKO؁�@C�2pڬ6�BX�и�7?7���N]-J�\�řg.��E��^}T0�@3=�B���s��kV�gXf�W�N��O����n���p��WTI&;2���ޜ�I;:�;����UnD�C;K�p�f�Vzm�r��K�ӟ��}c��O��*��dJ����)lLj��c�b��k��㮂Y�R-۱&V�ݑ�bR�'����$0������7+�1��`����bǀ�4E���v����G|�P�ܯ�9M��)�c�Ą����Abx�=�fD�7� ���gƂ�xz�J�݉��r�*�:;;��=�ǱWa9�@`�W�='�=f4d>�\{�\����1��(�:먪�ƍ+u	tD��tg��"#�B�w3*fB`D���-��O+���=��7���~���v�77f[�u |�/�%~؇�w���y�X$1��g�#�"�
��G�&���S���O� �hڊ((Q���T&!+��Й]�Z�ڙcDf ��8�hJ���ݛb5zh�hmZ��[�[g�߸�E���P��!Q]1�5�V�~���*��ۺ`��P��u�*[�+
����;i�6�sЀ��#4.�AB�+�l��Y�z��}��,`�~�I
J2�W�|�)�>5W7гsaʖh}h�%m��%tư�/½���01ȁ`~g�(岦y��������0ϱ�8��ZO�7b�G�L C>���3��N ��6��"������>B�@;x�=p���ş�tb�ɪ�yye�����*ȧ���\�35��?2ުfW�D��4�CFz��vt���^�����2��"T�5��
˂�8�"�j`s��v��7L5)��5�<�e���r5�k��������r�1+g��_���5�V��+�"��ӆ&�t���uK��Q�>
��y�������9���I��D�*@ǅ�0�=��*(�U(�{�F(ݵ��ˌH�=����hgqN���(s==���������4��\XZ���;)��|^z�5��ۗ�`/�K/��E���*ZW'�C\Dw�h@{`�es���A�/��3�y �Ź2�t��[���5>\�"�q����ٹ(��G�CY�A�4X�@�
���7�H�&���E�H~$��B�̵U�k>)�oO݅�����:�7��o�Ű�����}��ol}��ZJ���V��b�J�G�p.��F�Ӝ4�3�C���gy�
����!l�KQ6�-#7 �,W=�����A���췸�0��Y ��
K��F,���՟�������:Y�ΊUeja������=��Z��k��� �9�2x3��Y��j���2�&�xj�����W09�L�M'�r�jpC�����I`j�X(bN8��v�R��5�л����ҿ����w���JA����1�x���(H/RҞ���Ex1��7�G �*�Ot,��H���Y\�Ӊ!0�e��{���ļ����O�2s�d�%^ΪcD5��{��&�xu�E���k���lJV������}�"�
����E�#
͠�z<u �ʯ���Ѧ�����<+��!�X+���B��Y�
۔���	�Ko��(Q7x;,2��T0��c��/\���A�2�)�,��X0�A���/  S�f�*�������M]�������u�.��.Q����]��q��1��:�T��dʆ̀� �@�!a�ہP���w��Y�ۻ�g|�U vI<�W�lV�s��׀3�p�b�\IMך؟k7�>��f�B�T�'���j�7L�<ˠm@$�h�������c�#�g��m�Z��N�o��}�%���y���xa8���r��]m�.��M$ˈ��/�`�(���	�eKש�ϕ4@��\���8��F��:��"���u�����F��%�ei��ޗ��sR����a.��s��a]U��+.P@X���&���!�C��jB^`����I�d-�P
��O#V��,�t��w|�Q>�=.]�S�ص��%��Ӭ��v�q�������`r�M��)���<.�hlN/�#{`�JG-�A)9Ī1%��]��І(	:I�˰�Bvd�0�0��;�κN	��0-�M��3O�����@�����$��:����-�� P����P��K��h���^K:�A
�C�@1:�R*�fR?��v=�z�:���6�q9�_��͵Ⱦ��(�^��.U�d���� �im�!&�ĭG���\��OXA��S����9�o��a{|�j�g-�ݴ�Į	���Wg�#����e�w��vG끅�1_���j�X��V}�R�^|"Ѕ�����F��Kc��˗C}�0����G����ʌ�b�U�0>�j�\���NO�˜���c6-�:�6#�)��I��xr/S�n�|��V�=�o�����?��|=R1ٙ���n�U8���%T�eK�ʆ�;�~s�~��Ɯ�U������Q�JF��⩣��W)_1=�j'4�
\�����@#efgU�@��b�5b 	�+']?��~,�i���X >:�k�ʫφ)K�43�؝kg1�R��&�������<�SW�;�@,s�	ۭ�]�ELW��]|�ؗֈ�������O�TL(ሻn+�"����v�~z?��̛=	rF�R��K8pC��G�N�aQ��Q�d:���H4��SK��ۧ��g���F���	���0�������.�[TW�ɻ��ɷ}ձJ��Ho142�4��ѻI ��W��->��Q~��J2�F�Kx�Y�ƚ�R9S27��}��v��L/]�࢞K?y�rB܉���Q�3��p:{��% /��fϤs��W�>|Iޒ��.���Xu��~�DfK$ 0���X�c��qP5�[��ދc`N�p��bB�C���*fּa����dw�)L_��&�m|q!�}�¤T��\A���Nf���dr�;e�d��7�4MT.��Yl��]�^0W)aW���;�=w�Z����()�XJ׍����+~u��N
�9�MkaǹM�Ǿ������ڞy{b{b�r�&l��|���h@ޗ���������0����
�O|���XR��؊Џ��������,6��ƾ4J|�ޑM1�fU�ǚ��b�FYۧp��_�&��ˬE!�B��/������mǩ��u  ��غ��|�T��q)s�z7��\i^'��U_C�ٔ��7m���I}�=��a1VB�1��j_p]܀Q���{��$�/DF�G�l�k�.��Ȗʦ�t��R��\\59�/3���'����R�b��}kDrC(�b�H�i���U/+��Q�:,$��+��?��m�(�of�����_،޷�~C[��^��ֽ�m�Ro0I���G�L���Ru�����G�ؙ��tg	��&��,��%�z�;�.��tE9�	}(����t��P��� G}jjY�(�'��n��V|7�bۃ�|%��O�`��޾�-*�=Z�=2�ݠO��������������j�@'x�4����A�%�	�b�2���G������w_Y���Mw1���ݷ$)�@��  ��ЏM�76����K�\q1p���Ll<b���Te��R |sp�_'�=pg��9����`�,������~���� �)�'a��>�bC�!f�A��܊a]�8�=�7 �z/��L��A�B=b?��琱�'�
"��G�!~��)�j��)k�}���y3Ԫ�0�%�ǞS!��wX[8�a\G֋ǀA|A�*r�����}F+m�Е�Gr{r�
S�MV|��G"`%�J-)fo�bu�����][f�8>�_DG$ �r�3eZ���2l��G��aD*�f�Y��Y�"&���eH�?7�ss��h��J��v5�b�Z�O�F�:Z:o\�8p�ފ�����Ksĕw|�,����"�&� W�vo����)�)#��Q
����ш����sXU�ʖM IQ!¯R�Z7t��������Q!��P2Z��~���]=��ÀY��{�`��b��K[��R<���I����&MQ^_��j���0��kQ�RK�1>���
S�~*�� �[���0�=
ZƼLR����9*PY;�~����E`���<�����qV؃Y�~�_ n��z�>P�5
���Kѥ`1��-̸���|��
���#��OU$D7�L�+�d��9��N�^�B���d�i)l�d��p�����O���]���3�t��ġ���(io�N�E�#2R
�)uD[b�I�m'0	��]O1��u����~S}1>;���wR%X�`�C1�A�Z�\���vHFD���?y�)�J�!dkt�5nt󭋨�����w����0U���LqZ����df7Mw�?Ǖ�����^��ӫ0�Ӝ�����W$.G�v�4Z���A%y_�_��;h�.G��c�M�/����hJN�4�p����)��;{ h�s�@��K�����h��A=�J�|#?zib�رl��.�������~��6oƮ��r��ߣ�OD�0+fg����K`s���L1X���<Ĵlk�N��z�)ۢ�:8J��}��K�v +�;JXh&)3=��4�̂D�C�*�ЬCpgaK(�U()lW�X��hq�+:AN`-�]v����Ǯ�Iht�Q!��:ox5�/���,��ϴ�X�Z��Y� �_x�e�%w��O����oa�I+�e���G{�̶�:� #sR�>o��N���/����߹��F`4	ˉ�y���k���}��M��ypX�[<t�B�^�����0�!���p�B�ۤϋ8���ߍ���8q$J�3��DU��5��A��=u��ya;Һ�>�<�xإ���~v���ۖ<ԉN��6�ҏ�.F#
@]�d.�PB����p@uh��<���܏`k�2���SvV�� ��2�����&I	�=ϴ��t9Fݮj}K��D�|u$a�m����$λ�K�"�A����10���5���W��;{Q�LΒw6�Ѝ�h��u�Tc6���$�0�$�K8N�2��}�d�}��w�i�'S�^❩I�Ym���0d�)��Y�E y0�<ZjY��{;���$M��xX���{nU���<��@��4B�i�{��ߤVX�7]�4�_�:P����Ki��B�k���an�=�������8�K��\�1Pt��Ž��T��9��#��I�����K\�k��ʩfq��Q�K%��vv��q/���� � �@��v��t��ZE��d,@�0wZ�����<ge7��+\�F7|�E�3}y�����T�,���jn��٣�0���z�ɪ�~��dyW�k���m���(>�R:y��&8m�,Fq�&���_��@���U1��J�_�?�����	�9E�Ϯ����)��׳��`'�i/E�@n#�47s�Y;��.���R*�f��CXs���f$瓷 c�@M��YbS����7;�:���K`!a		J�ak��$T�u�>�ĉ0�d�޷r�����K��=��.���oL�>��@�������AU�	p�T��;��I,����G���x�.���%;1�5S�� -$:H�?�s'V������&&f�=k�$
��ֻL�4�:���*ҡ�F ��<���lS�sM���1���3Ӗ�l�����S';�_>������J���_(]�:ꜧ@W� 31c�q��v�M�Rn�]�ƚd��d<p|���SB�X�sL�<>la��-�p�;�b�� I��g9L�~��Ί%׹-��@�N�h�M�l��Q\g{�H�ߞgJ��5ƞ�1\��Ii�T;@�⌸���A��-e�Q�����_�&�Y%�N�˿^�,��?/>26�=w\�����1T��O��JV�����1��,���)��:T�����O	���</�l3��+���a`��`f�no<f� �	[`)P�n�iȻ�0��4K}��� �l���������0�n�m*$\����SJ��o�o	7-��\�J�.�+�6� G�-_h��Y9^��5G�Si��O$�*���u33�?X�@̧J,+~�{>P%J*l��H��K��(Nw���8��An~�y�|ՠ�dIr�XȦ�1�������4�~{V�~�QɕN�.ě��2��b�����l�.;��(�P6��%l��� t��Ϻ�jr#��wͧp@�� ��jDf�����t=�ٜ,�m��u�L��o�C�6�u�)�C"N�d\�i������JV�F:< DF��DZM6�^�9��}���Xb�m�ֽ*#��3t�a��������>:z�}�� -v,�x1��!8��3_��cǯ��.e��W�#�J�n�DxC�+��Jʍ��,����i��$eYU<u"^��ɳ�X�Ǒ��؏�r"/���D	
�vԈ�X7�Y.H4k�r���(`V��
�ʐԴ�	R��WSv-�S��{�z��/!��۫[�[2�e����X۶�/���(�Z\�z�繠h ��L��4��6N�-��D��J����;C���hټ�_�Y��|;\��
�������0ٲ�=���� �D�8��X��8C���8���7M�@�y�6Vb����4�Y���߈,WO.�'Ӫ_�eUb{3����[:�ҕ�y��.��oL[Þ�P�q�f�oݽZu���r#���ɞ�9)�!�v/D-�	�������yD tpf=�^����t��xC)�dO�Β�x�f㱆��v�e��e���	�~
���A��#/-�SB�Ɍ�^�x�{	�C$Gg"�_�t qR�O5����Q�)�Ug8��=<I��b|6h���b�Ԩ����	������'�n�r�ݶX���r�ۅ�%'�w�J
��9�H���1*2�/��''��ktDy�Z�~7��86��d/�^�!�P���Sǰ39v���s�H�	�� $�������C*����}G;���Zu��=��S��4�U?�̤����$vce�5�ȒG���L�����<�5?3t��A����TR<�숌T�g(�?�����;z�5���7�� &���a�-؆�pz�q=F�� o�=��s��aA�o
;��f#"��0�qd,+��Kw�5���G�1T���1$�~E�B̭�6M�
k�|������-�Q�E7)V���}���T�����Tٱ��&d���
S�V���G��U��
-�{�gz[%�&��)K�su�O�j>���<����	���$������$�����Vz ��<��Ǌ��>��}��쑅*։Jv�bc�~�4���^����g�2-ea�*�vzu�M��% �>\��V���
�Q��܇P:�lh^�=���_��*0�h�*�[�c�|�E0�#0}u��D_Q���Ye�"4���@��{�L@4d���*Aa�q�3>&��>άI�����2qr��=9�!�����g��������W`z���n��W���ܳ�T����PWfEtAP�2��y�ͺ`��F&�T-�*�?���������{iN*�w��⊲tÐ:���/�cNe��EB��N�,��K��8�cg�/U�ϣ��uk�4��%`e7|"ޭ��}����u5:��w/�>=�.P:WLN�N��`�>sJ�dD�Vi=XDvS(�Z]��|'9��\�,P�� ����Q&�л�(�5,������"tM��� ��Q�y�/v4��sy��lF��O��Ud �د峀5��@J��ڥ���8es@=_��ؘ	A@	���9�-!�U�U��DA1�o6S-?�h�M0(��n�-1��j3t�ތ�\���V������Ɔ������3��u\`	��#�������E����foI	,���M�/�m̟�#M0�%o�<�l}z*nR�њ2�\z�3m�ue�dX��6�K�E����| SaI���]F���3�Я N'y����9�
����Ǿ�p~�R�;��>953�;�I���dE�x_�P� �]N�T�������ʂ�M�X_�k�}���C����_�{0�h{6�R�%������4�(ᕜ��{�� ���}��%bh�$���ұg�_d����Gz}�xo�sq����(�{��f
�^�Ζm4(�I����������A�QI_}>�"��E�s�Y-�ǠI@6�[kwʻfaJ6����=�X%20!u�e�� ߑL��3I��5�D�-�X~:�n����Z*VT����j�@/�{0
Q ��3M�m~X�3�z��͍�E�_�� I6|������)�n��Č-B(��4����]���b��?��_����I����J�2쟲��}2n�A�>51&-��CP��p�����a`�K ��� n��"��?�`W�������x��_�G7e�	����<���x��n��)�OZ�ᶔ:��/1C���Z����*�k���/؈�d޺��R���X�[ʺ�Mh���%Α3�e*+Ǉ�<I>�0nz���:��[�0#I�[��?��7W��Z��(�w��P���b�tب���&���s*Dx0{�n|@�[U�V�Z�R���gvN�$%� ҙ�1$M��8���2]y셏K.qp8Z]�gMpPݵ^���89E�K�ZQ�h0�_)�:uJi�|�s�*ƈTc^��"�,}(K�^h#���ޭ�p+3my�I
��}�ZG�S���9?�Cx_��xE?��(y%�EoHe�R�P�BKA�o�yοO$�}�͝Buc8JK ���!ľ.Ҕ��֖	Ep߾r�%����[U�;A�yH�Z�{7�_󋾾��+��=��^���.^{1����b��{����R��tcH*��R�/Ѵ�'���|���opJ����3Gp�r�+�E&������� ���/�j`T�9��C�26<��Y=-gL�i����!�b�����C��DTɧ�`�8WW!%�P������,�/�X����$��%*c�m��W ����>=��1J��ij��y݌O��%���bTϚO�ô������Zأ����it���tq�������i�GhK�TU<sa�`~,�}��8����m�o���ā����\-��L�6$=W����)�0��V`��&��8��&�(�	�Ɲ+�����"���)��B�ϡ� �4�{�A�',u֔�qc�@զ@��:3��5�k�f�,��1�L_�5�DQ�ᪧ�f96� �w����uΈ�u\�'��ߴ�<�Q]܇ZX!ʤv~����Q����A^�aa�U;�MH=`��0ӻ�m�AI�&��T�AZͅЛZ6<s.U���=�1L�aaVZ����Lz�����9�B��H� mN�rnά�F.�sI��<E�� �Z����5��gR�oL������#B/⶯GT7b,l$c\?j����N3ov�y<���K�۱�ۛ��TX������n�:���ר"9)���t7�o��=�u��z��}4�_P{j�N,W�Sg�LL?!�C:� � IW�v�o��t��e^L���a��e���C����hp��SN%��PP��u͓�죄T�%�䯐~���p�`V�G�CJ������=ς�@�j�	����M9?~_�#k�G�>���H�w -H�G?O�[����?%�Y�笣��?k�5�~�d��]F�Т/ӽU/+������jk^�n	H[@ߛ��7����@ro�9S5ecJR �[�Vx��j����e���\�2��lTA��ߑ��S���p���>��cU��kw����P����eXf��6{	G�/Wd�SF���|�%�;'C��S�R�f6����x��,JA�~*^4�EVr�v�h�����������Q)�RjM5'���\�U�z�� ��$��iq`
f3w׈�m�n�]W`��,��.���~�(�?0�b�ы��Ø�l�
z,Sht.{�$�����f�	���|9��.5���F�ҖL�p«S-�����q���w|S齎���w�exL��J�Q`�� �[��l1@�pTr�"Z)�'{��_�X9��o���B>�q1At�?�,EݧF�%f�K{x����o�M�G��ӎDK���a<N�y�;����1<�^�3U���.�%9��=h��Ӥ�Z�]֩���R|�Y]������I!�`���"�E�-��Uw�=�5��F�	G,WD'[R�,A���|�ފd�f6][�^q������'����Y)-��ڂO�}�6���0����lG��n�b����6q+����*:j��+�CT�A�K�&G�hJn\�|k�%O��`k&��Y��]�/Sʺ2y��T/3!�L�����C�踩p@ν���J%���bpQ0�'W���[��,��A�H`�>c����p�9r(��{lM���"K-�6��+E�̙ݠ'q�R�ހ��wӲxV�0�&V�a�YŨzw5�g�8m~���On\����!bW+�:}q��]��흓Þ���?lI�l�|�PuG{�����h��7�,2���]dȾˍ�@�L��o�M��[�o�R�;���:�J�����}�2���3�Ȃ��]�v-�_��Hx�I?�ᾊ���Td[_�l7���H�1��d�nO�Px�j�ףqZ�����t�e����($"��-�>������Oqf,쿓�Ŀ����jَ�[�֬�͏	�Q��v]�⎼ne���M���M;�RQv$R�e�Ä�����Լ�2#�,�����M�cߵK�0���ͣ(���N�d�8%�Ԍ����.�$~M�Up��SHz��`7f��G�����9>��������f��-Ew^���ĉ7����.TT�_�Ҍa?�!ә�a"���9уs�G�m���yé�e�ձb��r/H���+��W��I'6$�0��i�_�9I�n'~�z�;}�է����~��^˻v������e�iN����c�����Bd*�T?���OA��aɡ�_�T&�ML��婸G���sv����r���̶��E��QD�Q�t��d��Z�z�^!,�1���e9Ξ��֯6ܧ ��~=@��Ph�#��3Q��F��N]�?i�<J��c;��ߩJ�@D4k=
`�|���F�(���|}��޼�^��<�m?���Q{����H�{Xx���I�	k��װ[W?�NUx�f�ȹ�g�ȃ��|t��|�yA�G����;���.�����L]g@SK�zp�WT�#]����H�%@�*R�HU��T��� ���*]BQB�Є�B�s�����_����g�yf��l�5�ʟU�����&IN�Ck�����~r�}EkĎ?/n�SU�����荗����X��7���[w"p���JzL;�^�"���ފ�j��`I�;��z���R����(S[Hș�Wӱv�xq��*K:k���#�1/ialU?���3����	���C\�d�򡶹>��\I5Ë:��Zx�bП�x-�#C�τE��:�E;A��A��!*��Rj��2��H%��/���,���%M�f&�:g?�,�B�F�CD�1Ĳ��oNm���h=Gm��f�Xv���S�0�Deݭ��P5��.�ZC���0�5���ӟW�pդ��E`���\�`�+����[�_L�/W��s4�u�p%�tj���ꃡ��<�aL�L�8m�����������<���Ǔ��,�¡չ=К>�(շ$�����F'�<CG����`ӛ��_�����|��%���ak0�X&6|�a��ҀxQc�𔲋�/d\�j�S�K#)h%�le��[-8��s;�^`%���9D���w�hzuJvP��UX���vJ���{j����w�{��?���,���w?�ΆPY���w�[ pgW/�F�à�&|��c�h��{�J�*N2q�JR}p��OwkON�S�����|%�c�_9�5�ܘ��-�㿙7q�H�L�G:���'U1i�C�x<�Y�����i��n���w� ��V�z�Q0j�����9�����C���Y�z"4D1Kv�x�8�b:�;Ow"o=�ey�ѬL����2���������v�,��q5W0G"��,�c�,H~���Y�=c��^������Z��Y�ŽmG�[�IX*�y+����N�k�2E�2C	R���b�������"BjI��+P��O��v�d��F[�����/�Q�N6�BO(���p�j�q����TNI�De{|��]�q�	����_dw��/����[��m����d.������d���W�G��
�� Ȼ�k��/��Rv��~�����p�1����PA��'O�Y���`�Ef��ӧ��^��3�^����ͲK�oM�@5��im%4�C��٫0��T?W!()	j,iF`:�dW��aQ/���k�S���R�����S�/�:Q��z�~��_ӘO��hN�B����w�臒/�3(��%�]���}������l�;S����6�#��OR�2���)Kfd$�[����Ǝ�M8��)Rᡄ?�*[L�$'�tL�-��d���$�oX  =��w��7���Y���jK��qP{�s��h�R�ehȍ�w�q 	ժ1ۅ���rL�.o:�դ)[*�P��QO%�`��O��HH �F�ͤe5�Q�p/���b3	���EHL�#n�{.��FD�do۹?�j�����<$2�CO���kE*�~�����Y��Crá���/M�k�gቢ��/:ܥ��82�I=q�ܨ�#���my��Q�~S�\2(��`:��p� �wH����UR��j�nOB�CO5��[K�\5}��6^�ýt��Gv2U�=��rM��mԺ��K��ˎ�rF_|��Jz��bה�,ڹI��ڷEY8s��˗]̤w>�b�@��r�H/j�iLY������&�r������l�ܝH1n�R�~;
״���KL�Qo]e�[TVx���Z�3�l�V�����2U�
��g����I���:�w�4ńN���;*��.1�>4��{�LLf�잦|��7�|8ו�*��X�qys����F<�n��@A�M�0g����p���j��c��֛�N��}�'
y!r��ñ�x�4a�RH���5�<���kQ�i��]a;�ұ�ר�zxv���G��\���0�J5�!��Gn1\[�{Wlne� �ֈ63力������:�j�A��,��nZ4��:B��!��~�s��E6��~���k9���q���)�uAuQ�Bߴ�w��s�}�'�'���1S\�����t�s×r���IGs�!?�o��n_Mk��l$<�YX#q��F,��V'�gT�O'3������홚S'��u�:�o[xڂ�֪�nb��+$3������G/��y_3�|a�[TS��^͕l�<m ګ�Ng݅�-��b��ܧ�aGX+B|�``��dm4��^p�.b�o��B��S5��B=��C�4�J~�_ۚ�",���th����]�$�v��c���n�P8d��?7���`��r	�R[�;E*f�M�F�R���e�M�����K�\j����/�����9 ��)h���r��T�����.$�4�nLn��¹�����*1��?����s��e��{eQ��S��l�����|����,!�:�{�~o!�J�e�Ulg�FV�>Io��0�W3��9Xp���ҽ�m����(�^&E]��-�*�{���4��nǔJ1S���
6����8΃�߇B|B��T~�@_D�a%o�������exa�����.D|�(�r��Q	�~���~�z��0������@�?T̀�t��i�.��x�2,)����q�6�~V��:�g�S�+�J`U����������B��I��Q�;/�wj	����*� ��̝�.�f�c���'����졧����K=��/���'~�͝:ع�͌������Oy��8�����H�!)|�{�uS���$�t;-�:����.�X?�=�,^Xmdˏ"�=���y���j<G���A0�<��d8����������#��MUbp� �irgP�Wv&���_�Ty{����Ub�a Csc�
�mK�F�"������lV�(���X?���f�e�j]#�c�}a�k`3� S��%��T{7��z{������j;)��&�[u@�ؘA���܏ˑu5R���<-}� l߻��(^�tW6�&,�*����{��R�ù��g�����&�k�Hy%y@v9S׹�+�X��]!�rݗ"�Dn�ٔ,尞��.�T�v�j���9f� R-{�폿F����"���h�rs��5��{�$��6{��🙏�<>z���i���&7g������z���$�2z�V�a\�i�_"����^�D��!�=p$#Ƽ#�Y�5�;�ʥu�DR���3��\y�Nuk"��J���ߔ�b]��	������� U�:�ͺ� �OR�FKLב�2�{(S��)���,�6��4�Epq2Q�����ґM��&yl]� �9�F�a�ȥ���8�d����>�:���=�9�5��R�nkF&�i竷?b(�4n�IM����FU&��'��Jz��E�{ y�6���7�L~��[d�0'��tXVb`���(���Q8/�����K�Y���b��6J��6a�C�в.aN0l(����0��F$%��)w��4A�C!"
��g�ٱQ]�j��O:ʮR��SZ���(��j��<�����M9�]m94�!rlA��U����M�YC�Ő�N�ڊR�d)�j����BOdꩄ�����y�wI�/�A?0�暆x��j)�~�F��K��r׍���w.,�P<靬��������� ���l}����#�2�u�x��;t�T�@پS�q�q����A�܁Ef��|���l�׀Ph.��h�\��F�g�۫.�r&a������-r�\X����t�0M�iD�v�@�*�|y	��]�MO8?^�H辐�6&(.\OpM��e&���0}��L9n�F�j�����Zy��(?��!iy�g*��u��]��A�H!�{�d�};L����'��_��6�|�z�#�R#�C'�ö��F��&"�+Q�&^��@�I��1P>��N���2n`0�Nh�q�8�A[Š��9,*rf#��3,C� Ȟ]UW<~������j��hZ�����)�)Z��+ǜ�����閕�����
�J- ����m�a]&&�*)��^��g.�5�S�(�uR��y=�3����Wz��Op��LR*]
�F4X	8�᡽[�Cjʳ.#�A����Jg�f�|8���m���`$���\����Մ��/@(��髊��B{�81��,eg:ږ��^ؓk�����)>½qw_qcLy�7ִ�����*�F+�_�Nz$���%P�bܡ�mQh�{�QH1L�Kr��G.;JVPP�ӻ7�d?nw����)���G쎢��:��8q[ա��@���##t�~((5��Zb���g�=�]
���:!T.ܨf|~����["e����L3_��s�=�$=E7&��m��w������4]�wvDu�Q�Qo����(wJg�a�'MS��rW|h��?���ri>!���#���U��j�k�.���x��ZW1`�9y�x?��Iʩ����yR��g���P� 
̋��5����/ov��+X�Fp���^��؀��=�T]נ����)��T��.0
v�����L�)�Jn_S�hn:S�(}���eV7�J�F�uj��;����kzG���nρ�����g#��{�pW���������("��S�n�O��r#��0�� mM��
����<g*\2�Cʪ��t���1̸RQt|p�DT�����9�.����l���2�m�{�4"C^^uN�j��� z-�mexlnC�,Ě�mM�	�2~%t@}�#T���1ԕ�� ��2%��v�>hD{��m���9����0})*���ٸEr�ۯ�_w���lqj��L`�2�#���7�����8�Zbo��!�"�lI�Q������p9�f���z�h�:�3T:^�%i���CL���V��I�f �����
 ?�V� ���ٯ��������"j�J�j�1`�+OU]�	���&��$���o� �>�r��ӫ��:T0����{�q�[!A����P�S��B_5��	�.\.x-�,��&�cQA�۩<ˏ�D�t�����x�}�;Y,��s��,�&y�_���2��`_���������0ec@����U���)��az��ś��DG����z�@?��n�ݬ� �*1c`����|���U=]����>�z$ʏ8D�O����1�L�Y��pTh�s�؞vL�z��2���Ӳ�,8������ah��z;���������rz���e�$ߧD?�z�qAXJU2�4�xSx����ԣZ[,v_�E<���A|�T �*m:^�p��B�+<�]NԵ$�E%����1fU�1!�8ꦵ RWQF�P@���['�z�{����L\�g�Pu��r�MExkOB����aJ�xi35˒�D��&%�Q>o��]����j��r�vmI���-{�tN��_i��.p�c�*IN�(v��=�K��4���{1�� ~� ���N�MNޱ��֡��,yv�o�%�<땘eQ�n��Aj���E%���:_�t[�|l������ش&�m=KrI]"�J2���v.����/B5�>�����D:�*�ѵ����cB�3��j��
-�md���F�w��SAv/�D��y`�X�BST����H{���y���G.�:z�r�Ʒ{�[q
�g<7�N8�r��V�����?_��=	��aJϺ*C_�k�J���2�O�	������N��w ������_V�ߌ3z��#Ǥ&��T{����[;�q��do��M��nRC�@���i�U���&����>k7�\pB�>���	?r#3͇'N��!�g8�S�2�+�;�h޵�M�.�1㹕z����% F���V���F��Kn��H�<�*�����.{K/jq;Jͤ�Zp��I�`�}��3�/�veZx��g�� ��XL(��	g�P}�/�?$u�KWn�x�neMyG�6���j7<��C��i�n�:TmE�y�
�"�����Y�DR~/����	쓜�7ZN���ݪ�u�_�A�+<m#	.W�*��[U���k�/#?����|E n�������P&8}ڴ���١^�T-��_�CC�'5�(�������8r.����p���0h=���"W?��九92j�Q	�`#8��j��:&4J�^]�Lv�ڮ"�^`2�}YnKy�`����j�����,3�f{�+���\�"2n�^(��}M���΢�}�ۀ��8��p����
�Qe`5m�������M�򑬲�	�K+�����%H��q�É�����,�X�K�7�lPsç�څY�
%K���K7�����r���k�5�|���������X�>s�V��m�&2i��Y�>f���j�[M�QS�����ޠ.H�ʻ��[ėԺ�c�D�2�[��F�MI�4[��G�ؤ�
e^k���'�H�)M�1h3��YL!�J~d��#���i�hu���l��GF$��|��]U�(�4h�2��ת�:����P]cW����9��3���N�QI�G�L�dW'����˛�C#���N�\v��O\�?9���_���¸FX���Ϭ%�]��g���eO�a���	YJC�Т8ز!@�Zʟ�,�HK�	>�nJ<��$������y�W�`M�HSf<���a#���gx��P�^$�~6�-(74��FI1y3Ћ�gc9������+]�-�0W0�F$wΠJ��� ����e�N���|Q��m�]�jS��$
���C����j�2����/9�G���i�z77�J3�|I��̘��KD�����*����#��d����1�c��M�6nfk��y:|�f�慽���{G���lYa¼�9����痍��e����A�nGnj���G�\YS
����r�˸���������z�|���PY��~L�,[�u�Ӎ��z��2)4���}�c�7���"#u��4(XD����W�gs��Ն��Y�渽_���T�1�(�,�M�u��n������9 #���,�����Z�3���FB���o��IĬ8�dx��e�]�ɗ�.����Ӹqw�:�j��DͷM�gHс!^rݠj��W*���RTf�G_.k�qs�P�rØ�5���W*��,�}߷��%~ ����;��u3�9yJ~^}�ߨP����1��*�%[�6d�q�ɼ88�}���l�@,p�qP��l�;L�C�Y6���������C�{9�����oR3)���v�������l�_Բ�z�6����>�Qg��;0�6*R��P$q�CTJ(�W�iŐ�>n	�#T�O�0}3ں����0�=������5:�y@�d�&P� �ƻT��)�R5䗖�r���X������U�Z�o�p�e-��z�ㄇ��J,�����N�Z$���a>�G>��?M+_a9��Ѥ��\ڼnĂ�-	�M���Ɨ�3��8��^,������v�R��f�/�W���C�F7��}Ɨ���Mi�
)�ZZC�}��(�C��eٵ*_��~�oOIs?�Q�k:��f�!��b��^�d�Y�x�AQd�2�\�	�K�1|�,<'&�IPG��{���c9�o�Nyp���pA6��國�rp}o�ދA��ܢ�-��z�;�d�*�� 8)�Ƃ\
I��[&��ܬ:3D�E�lne�i�ť�]5�18۵��L#?��6��f��t+ �E����*���"���b����?�e�!��3��v0������0���nￛ"U��X���6���l���E�h� �b��4�c�>q�R�#ұ�g��Mr�:,9K� W�(n%,P�U�ۭkO[6C��vEwx�����K�)�k�^��:�fB�D��[$hKM��m���L�d	���\��u�gX�(�Pi!�d�������T�3BnrM��4n0�n�.w�[e��c�G�긆_�Ҿ���I|�;w3��rQwb��ln��0_��@��Y�Qu�o�x����<3�����R2�aBh��X��ݖEn2���(�epdT0��(�.:�A�˲�_�}�4-��P�	[��"�R�@Y�=?ˇ���L����d��G�tϘ��B�kD�|�J�1)�]?�k���T(1�8r���͘�[_�姧Y�J��o�w��� )ȕkn����+��)Ϳ���+DV.2Ⱥ��od����I���G�o��MQ�oˢ��8��1�JJ@���==fQ�����+�\	�x��gW$}M�V�'+n��2 ��ضi_�?�j@��1;Q�e~�,�=�vX����Dc��+�!@�W�7́����]��GG�� o*�\�E��4 ^-�p��`�j��綛���g���Ik�kqN"!y*�۫������M�hXq3�������LU/y4ÂWsbb��3���""\�jo��T����<�?03�0�|�ċ޺L�q���ejw[�bej�0�f�|���mI�$s&���l-<x��Q����Q���f��\�ࢥ��^rrm�H����n�@�٣R0���U���I�?�S`Zn\/�vhls����xteed�3S�|ߺ�ұi��@,|1'\�2h�b����!n7�������O�P�ݫ�XZ�����Ր�Q�Uh��8 �[K�����WVG��ip��Y��ay˽
R�h�oX�� �Z�f��Hi�\,9� �"�Qt��9S �"�����BYt'c�ٴL"�DR<�J=�9z��P
]�/$mT��h�����w�7|=IN;�MXk�T�)ﺆ݃�f��.����7e�V���>�Z*A�l�=;ԩ�:|�=�����J�M^d��J��Zښ̴�s:=�5��p`���Ȱ�T�3�����%�O:�ԭ�o=2�o[�p��d�x�`�)]L�<G��	(R���v���)p];��4�4j)L�&ni�~I�5b��j�M�`����}���鞞^77�@-���Z��XN�u�Sƀ޵�=}�1�<��'�X��ĳ�~�D�1�-Z*C�$I^8��UT�^Z�?�eb�|�%�?}�4koi(h�K�pZ��ucHYz&�Z�ɮ�h
�"d[��=����'�@p��-���VA����ժ�����IC�����:6�g� ����v�*�i͚O�OK/�?@�Ȍ6s�jR�念\cֈ�si>�,m��ѓ�)5�����Y������Eù�=����{k��a�j(t�	���R��j��K6HWٴhZ�����9����}
�G>M�=Q�ӳ�q���y<�⡱�Yx��EFOq�N��	��n<�:��r��K>�Q=uܲ�(�Nr��I# �rD��R�i%���կ���UC��Eg<�
��@��H��"��Va�J���}᭐ІM�����<�&��2�H�ť-��n'��s��嗇�t��-�H�\:�1�(\7����ď�V�^|�%ZǑvN`�ʥ}��Y��Jwu`$�M��GH[�/5[hu�ʹ5��0P��m�� 0��t���e�ǐS휜�˸)\]��`˸�]Q�������/��h��i<b�'��vdAG���+��h�í���q���e�%��l^I?��H��r#N�+�`�w�W�TJ�T(�t ox�S|(��*���H	G�f<�蛉�ͣ@�6U�S�#��!�tX�q�B��S{E��mu�l��˧�&d��?V\���՜�_)�S>vr4=�'3���H�MԆ������j������z�M~��OSx�jy�֣�G��m��0��cy�XB��Ǹ^,>�l��I���E:y��rǙw�<����s��%�o�s<���ETiD^R�o/��Z��WF�7�	<�t{-2@��:�V��Ώ�5�["��a���6M�]����W;����}�rC��=��<���B����T�~뾢��+Ktg����³h�9����+$��\��!�2�S�w"�D��u�m�=�Ğ]��V�ĵ���cl�6t\2��A&+���< �[��f����6�@�����q3��q���!��߇��τ�.
B,���NdJx5�>�����s�9�i��C���v��l�0��3�۲rV�����!�l<x���隥�쐊6���=I�6��~Z�#�
OZ�'��2C˹���W$+���z:.ӮJ��!�>�W��𦸵ȟ��]�7;�r3v�9�f�ˬH��\�P�^��䰾�#�;�w��B���&n�������i=�q�V�}��"$Y͑O3�M��c;2<��\.�Q�3@J޻�:��m�.�:Bg���E��b����n�'���)�Ma}�Y_z+��:gW�~O	�����ًɿt� A�7ɘ͸:GH�L0�8�,�4���"�tzYr���V,\n���+ �D� -^J�4-�:�ݯj�*/̥��3��a��L���c8Mw�"�0����n0*��/�=3[��`����m�Q�@RL�����5���w�`jøn� ˓���t����t�뷘_Ѿ����ʼ�r��{���j+�٠��m�0g�2��|�w|xhP���FS��>�ҵ���i�["K yzP�&��q�=�����G?��yK�Y���)n����0C8����J��/{�� 'Ɍ:-\Y8�O ���N�B�
���sz����c3-�F���Ua\;oh���YeUO�f{�	&�O��ٶ��"��Sސ�ָ�{&�x�Ǜ�׽������9:-x&�;�V�k� ӓ���4QS4�rP�$�*ll(��IK��]?�R���ȓ��*�W�G=+�Wl6P]n[zl��J̔C]�=���*X{r��FjLaC�<�K��v�0�j�|4��|�K�����>�����m����J~�Di��f�!�P�q��3��5�T�
>��bJ
����W=�	��=q�8�7���6��K`��U�m�T�0�B��x�m���>V���@�CZ��2���f��+�)\˯n���|�f�_s����̳����@h`.�k�X����~j�/Q�5��&��c�������A?�4���e�|\���M߱�0�vN���2d$K\2#Xks}Jz�n(�$���d=p#=�I�i~.�yb#��v�w4��{`�3�tI"N*˒*5&��U�9��h�n��_�0	���� Pzu\�lWn/h�-�,����14�R^u�����q�h4��6mR{6�/ņa
�qkc���ר�r�(��y ��-%1˯4'];�4S��wJ���2K�l��@P���Az4f���H�)�  ��c��UP�c�%�V|fy�j��nn�^,n��bR����u�ྼ�*N�}4dEyU�_7�.��{O]�>݃�8��*>��Mw��?�J��kb�{�t9����� 5e�(i?(��:ވ���TmuB��Ƅ�����YՊ�6�_��tF��̯c��R,Ym9���{��O 6����t�	y\�ԧ!n���	��8�4����(�NA�\���y13�S"\�Rk�b�����Xu�:�e��k���Mײ+BQx�<�4Ģ����z��Ew>��?�����)�F��
Q��k��e\��$��d����F�ǢK�����v߳_�i�c�~o�.f�U�œ�Nf.����_���P
�%��v�<�v����4+&��V�v珙��̳츝��E)��@����r�c�V�*�7�p9�~���^�w��;x��6jH>��{���m�R.H�+����V`w &��2���7�u�o����1}�u/8K�4���۩�z�B���ӂ������6Q�<��u�#�M<(~,`�C1 �����T�c(�C|��2Tx�*�$~�:���؈|�R�~����^�{P�y �W�W���8OK���Z��v~9����^=�k�qmJ��,�_�
x�+@��X�zpSN�h�����N���v%�~�S_Z����l[07����	�ҹ�3��0�@�Х�zG���ZG^�s8H��s %�����G�Cr&�V�&-��9uvQ���.�w���e� ���5��-.٠u�+�)yx
��NC���c��FD�Ip����@4�����[�:\�-��� j������,S�c���"��Q��THK��{�2�[,ݾ6$��e�Oy�*�8>��5�a���V��S0��8q<��L<���"�3���Ȏ�=�����a;��ɷl0�@�!��1W=�nB�|�����y$�o�e�[�*��9
�ۓ���v�����D\��1A�(T���_C8��ǣnk�Q�����z�6 �n��%����c���E �f��o��[)�;�<ƠX�%�j�}�x��
�mWc��w����-��S[��Ϙp�H�.Xe��3�@�.��F�����HCc���*�n�Z�t�%.��᭣�Zya��ae��q�5]�$l�F��&��⨛�I,�E-��\�cbX����o���S���?�QN���Ժ�ks�FHRl�j���Y��a���+��<�z`�-�3j�ghy_��Q>+�PgQ��vI_��b�G�u>:�����W�9S'}��L;���u~��,t&:�Czh��A��?����龜����옸��EM��>P�U����	���%��6x�uN�c;@=�
F[��1��l����2��m,�����Zz��ޞ_n��J������߂���	j���NC�b:%3>��nH'<�z��_a�����n�J�������3��z�����NJ������v���a�V��!��(����N.�ܧR_@����ur�]K�Հ�N,��N/�i����C#�ZgL($)9RWH�le���z������'�����J�B���z�ݍ1p�N�c�����Y}ݣ���K+�xj-Q���� �)`3d^���LD���^{Ę�
Ÿ6�!~m������Pl����D��聕8$���<ӳ뒝�P�����C� -wo�p��� 1P��waq@PS��ߺǪ�-Z�e�{���:��=��ۀև���+\�1 R;i ���"6������"�/�!�WAB��؂û�����pk��<+��x����h�mI�+a_�6KG���͓����]m�bd��҃wL�4�
P�v�ߎ�M\?I۬�ߥ�����)��K�k&^c�om��$8���x��L���5$.P٬	�0����H���	_��/f3ҼU�+���	��	��ՖM��񣅹x.������Ā˩<Q�7�6�k�,��-m*������C�!Է�~�0��AsKDJ����!���֝�)��_�P?��_�����g7FH����}m�2�)�I,w���v��݇+^�˱C��9Zq^1zQ,-����)B�>��U����"D3�x��C����_�������m�S��K�������h�aQ���ߝ.�����s`wu��aٔI^V��r@��P�{hDw��ni��7C%��Vϵ7���f\z��� #}���&�*h�k%�o���kR�\��i�
c�i��)��Wzw>��2�AuXg����i)�B3�(���~��a���Dǳs�]��"�跎U<p$g��˃!��Ѿܳ�G�.�=Ui��@|�̜>i�tB�s���5J��l
_}���rE�&�Zh��'��	'o�E�I#C�;��;$��|wY��V�?��c�8=���My-ˋ��Ňb��r(�������
�2��2�����r����wg"�d��D�Z�<x^�W5����i�^�'�~��]�ܯ�a�-4gVn�k䪧)���4��[�4���
�m}:��O+��6N I�꒸zǑ����A:� ӕ���A�]��#{5��AU��������mA0q�ˑ"�Db[7f������L���gMĨ6� ��	>�&����	d�'j�G�P�Y�uŞ9�X0���LjP��O�`F�#-��9���ZOB��]��qχQW�a�h�>%�w�x����0�?]��B��NB׳2�jeo|fWج��$m�zL8�8���傹�]��'�ý��|���{��~	�3��9q�sH^��1D)�	�b_V/�5��{�L/�B��O���u�����	�a��D|�ޱǉ�[UW����.=3������YY�֨��D
r7��߁�__a%cup�(�?Q���v����%�5�v�[5�VR�%���w���]�����������g�Z��r������B����Qz'�g�gәF����&k������[��+������+�NV8�%�+8;R��h�>�ޢ=m�KK����Jĸ��Z�.BJ%��U�vj/��^�Ul���s8G����ܦ3�c��@�^/:-\��k5�{.��C��rʩ�֬�/���ؓ�������(��{�����L#�WLe��o��#��3�Qc��Ӕ�$|3����Ck�ˏ�z��woGu/�{�͉@XB���חS��d�lr{u2�0.݀� ����#�=e���6�u��t�?��^r��ׅ.hOJ*��v�Q�a��!������\���Z���zr�=C�ϋ�8��J���L��$mK�	�M��u�Kq�
���r��?�/١+��V5��BOW!����u�!��=�j	"lҁ���`�/����)���Wf+�j}4��(,)怤zQ�;�a��� 6a��7R�"7�����z]`��gϦڥ2��#�K2��R8�,Hb�b~ 8�,��2k�+�ئ�ү����x}˒�����j���oy�h�j��\z�i���*�����+��I�<Qh�l�n,�q"�)�h�y�b+�~-v)X�v��(+&���U�މ$,z��˖�rM3gֲw�I/�
��NN����n��-%h]jah��L�.�rl�5�@\[��B�0���޳�?YvӘ3@��ϛ�1�=^c�w��O�~��Z6��H��	�]5�T ^�J�b9��o�0p��/{�!��R���Æ�:��9�����r%�h�_�2!C����.��aNw�o�8|P�,Q�-�W�����`�e��OU<��<zE �.����1�D��N������� N �:K�d-J���s�X�ǩY�R���<7�>>`~jݬ �;<C����߳��������@V�Cw�D�� �i�ɉuA���>�_pY����n0ѱ��dK���zg��|�G�gg�%������瀢:����C�h46��wPa�sML���.C��oQy�ޤ�lmBF�X��o�+��D���y���G�2Y |�k����w����"/8���`#z�1��E:?�.��]v-���ߔ���s��v���w4�<�eWg�?�OG����M�*D��	�	�X��n<uL�E7�eJ�0���L��̣E��]!7bQ{��D�@��k��)����u� ^!�J ��{`e�&�צjPHƄ`�� ���ek�Tr"c�Z:Y9p�������ο�D�|	BC���[mת�%�Q<l�.1�	���	��=jZ����� !����������p%V��Ȃ{2L�W� ����w @�e�0�Ճ'�  !����Hl� }%��V-Μ�K�dM��r�jxj]�Y��!�� ��a�y��}���<���{G�8�gN�����㗘��mA�oN���W�R>^V���c��Nʊ�v�Ʃ�W�� [��p�o[�9Xԝ�4d�$ߗ2;���K?�#U"?��É�h�& �!�3yh�t��'Jb�3�����r�3�]��� ƽW	?W���F�/���Dw���y�f����7�R��W�X�����V�i˦p��4�)5Z_\��O;`�n?��M8�2�#C��j�|'2�$�L�$A��/�\���hMkܛKe����9�>w���t:���PQ���Ć�9t�5�c��8��x4D��]���>Ϛ�SnepK�n� c�T2q�&RA�au����;㟚�wm�#냸��5�Q'D��/L����h�����G��c���j��<H^�����ۛ�D�,ub���v#PE�\�IN�� �C�?ﲨ�M��2���������Mg�z�j�'Qv�X�C�$��b2f�r�voX�P�q�x #:Y>����7*Ȝ�k��9�Z(g�k�,*��n�I�ټ�cT%+�8��$SߖbX{*�'n޽�p�, O��������W�h��I
5��cH�	�leo�Ff�>�����'� �M���e~P��G�2��1�I6���N���]6.5�s�Er���W�I�t�B�+�?�}�N�'�	R�<���go���;A���q&N��t�p�	.ţKHjhV6����S5��6Q6{=4� p.O��U�H�����J�>ݡ+���/�p�W��8_�žl������`�'�f���ζ�)�u]��A@]��Y� .+@�����q�Չˊ8F�V(��$��
P��=?�&��N�|��
=����ey��*��3��|��mrl�<ɝ�����9���N��J?����X�H�m�L�̬��l�/�)ܖ�nTÑ��+���ly��ﶤ��o4����oe}s��]O�9�ԧ��M��L���A�{jм87`v�U;qY�V�S��B��wN�
p�2��]-oD5}eUߺ�[��~W~H+�:A�i.����N�b5˺��Vf� ��X5�+?�U~�x�4Nw��[��Åμ���n^�I��0��-��^Sצ��?5�R���9@HH���2ܠ/:����K�=u߲�����ŰgZm�d؞��@Q\�@���
�v�I��[(F���@L�AC����z�J&�z�#-�f�<�U$���C���u]�������M|<O�@jLH��J�'��>S������U�$��N�?K�L��Y?�-�:x�<�^�` ���sb�H86$�`�=o�D��D,�����=t��S��[�3�x{1I�s^�.����Q��=QI�q���0=Π2O~ȃ�v;[2Yҳ�b׎ȀF�?'x&�EH:�<j<�:�u����0�8�L�G�ηؘ0V�=M��<�c�5^�C~S�G���v�_���+Z�����h�p�Ŗxg4\�r��~4%G؛�g��{���ng����m�I����i	h=�T��m�=ώCR�5�3q��!On��v衤l���]����W"�WC�E ̾��Z�=:������g��V�m��x��]��!���M��"�z$�!�qג�3u-����}�kC�va�=V�泽�Ь�,�����S/>�9zj��\��nGTd��4�?^������	�;�=�nri�ə��I㧐�S�Bu��(��[�?[WW0"��2A����I`��sһ'��H� ��svt=*[�W�V�)��(�[i���@E������~U�H�Ʀ���4���Q	Zƃ_�2(uّ�}����Zٶ�ƇP,�*���}-�-H��g�6��oL��DG;�W y3z]}X�Q�Au@��+[�E��Պ�'����.|`\F�ߧ<���gHI,]`�_5�&5T*	y.�`�@�pk�QC`�'���g��%`��	���y��*��Q5�Ŭ�O��"��\5�}�O�LZ���/��R�<Ǚ�����Y���&�����3S���QK�R.e#�u�ǽ��Dq���T,x�s���q11����f�]�K��Z4���}$��ɋdPd�	�}�`}�b-K�tW�o�w����H ��ߌw�֨`�(�9k�R�^N�����F�KRj�T�>�L���rn��F�g�q���ގD�O=j�TZ~3�3�="/����N�x5��������jj�@��("�T�"�;bA�Ҥ�*���(���B�J tE��4�I �5@���;��{o�;��u֚kι��guA���:
���[9ILay����Y�e��~�x���� �݀�B��lxE��
;\�tV0��|d����JF;,N#���#�k���?I<�\�72�5�+,�UX����lW�LKvҩ���*�eC��g���Tf ��Z���|����5�z����l8\Y$o��D��C7:��P����V�b�d.}�,�	/�啿�t8�����3` kTR��|>8�տ5��ok���~^@*-����{��P�n�km�}��*TM���>m��>��r�B����V��E]�\Q�����E@DX�
@ح�����U��^�sBo���� ��Ҥ�b��[F�L���0Li�9}�T�#�,Y�0��T*1�ߪ���S*����7G��Qe��*<�*�b8�� �7�4n+��dOU��	�QȾ�K��#�����초�J¢��t�����#3�K�b�j"R*/d�����<�_y{��%\K�`.&�*� �4c/VUA��B��U%����;�f�=g��1��fթ�ˠRl�␆�V�VG���v�� Iqm�r���y���W!"c�3��6����}V5����H�E��&�bbc��~�{���Mfz��3S2��qo�Y��rNf3Kvro�	�����em�!,;����f&н�>A���aM����(���}%ܨK^�hL8��'r�������i��
�m*��#�ި�xs
J>�b��џC�@�(`���*0C$���M�c�N��d�72櫵�o�/�ha�d$�������R��VX�*˜a�S�m1���i�%r�aV:����]y�f��op%��P����"�<P�͸�?P�>����kl��[7�&f�O����4c�����O�,r��wk�%.��$�eB�ŀ�'����O���7�{,��t7��fÝ�����Oob�|%p7��%���=[5�~��1&�i������A�?�X��!_+�'���Co��6̖ȷ6���o�B���^�6
��>�_��48L�`]u6j�4����>91M�D�I��M<�It�w]0k�j9rf�D��v*¥�DSlM��T9�E�}�I��(OY	�n�J�N5����q�7�'N%����0�Z���:�9r���+b�3x�D.��<����G��:7=t{���.ѹ��	��,���h��YҺ��,��&l���J�����r0��̮�N���"�>���Y6�x���i�ƙPAl���g�jA~�ĄK(�z5��'S,~a�ɢ��/[?Sizf"���ֺ\�<U�:�I<�cP��6:"����+�x^7�[�TafM���V��)����g��R6��#v2;�m1f�E����9������2�r�Na���?N_?�q�����݀V`�o�E�W�943�(���s�ns�Z��z>FB#/�efg�7���A(���Pb�X��.���K�÷�N�??H�"�����9�k����+Z�������ŘE:ঌ�y���G�$ۤ�ڋ]<Y�c���T�4��vP#��!�Ib{��Q۱�	�7��u7x�-u_i���q��9�4N���$`�E�ǟ��wZ�M�L�� ��1� #Py���b�М��Li�z���у�-j������[���5d[탵���ӥ5 ���w 3:�%?s��O��C�x�j�E����'~"�^Ti��H��7]<5����Җm'}m�=��N�,HU�2��*`o�Ԧ��:��Ur��hgw}��͍�!'F4qrnI2`��,���{CS,+W1!b�8��(*�	 �r�����6�x,c)sz�Q����>�,8X����f����Rk <�]po�����u;V�X?��S;���߯��� -t�g�?D�#pyIm*�14�W=�%����:��B�
�fꧢ�B�WO~��d�_1��:�CDe�$X�F(*�c	�)ڃ�,A�]�����RR^�6��䈟BO.�t�=)���'��H�Dj�eK}Ǧ!}\�YX�qq�K��̢:��30����x�
�䇻)/��$[o%��YV�w96�g����ES�os&~a���2�.9&�f���u��I����o���/�E���o��;�n0��D]�v��"G�'�ceKp����g� �\��Ԭ��}O�$����R�ud�Bo��m'��@Z��p>m�tI��:�/k\@����~����,�`��i��l�%�q&ދ�87黊>�)�5��G�!i�S��1h%��Ƴ�/�� ��dY��v�|�d7;\Us��l�����f%F>Ӕ1{	1���9�C]��mh��BqӲ�����7ַ�������(��@B��U�|���{�ؠ"뫺�TBj������WS#���3��Df���E'���O�f�N
1t�K�RG���G�t��6�O�V�L�o" q��q���0�Woѭ�{�D��k
W��Ơ��?RY��*�
;����>M�e��s�-�lc���s�1V��3~�̫��o�����r�"���N�i��q�����NoB�P+�Qof.�
`"Zش�?�w]X�eE���`D`��r)`������j��)V�/+���>t�>Qi��L���P���J4������)������12�[Z{n�	�B����;�K��"�<kۺ���\o	�f���� ��4=���q����o�=��<����j�S��	��}���̡M;��q�����]ٖX��Jgk��05I`ZykH�[�=��������ɭW��g�vb�	=K=�aq#����zY��G+�sù�1C���O#��t^b��j�	�����rBw��5��/�}:�X�Wl��E����J��\��Y��F4��Z�'V\%���y�J�L��W$�-���y����ܝL/2/g�5[�;���¥f;g�43�'�Y�̵�����ɎN�#�jR-|�-)o]��!�E�'��D��D�0���1��UҫR�XD�}e��68�����Hm�O �}��o�~{�L��l��✢�����-��i�T���cei)���[���?�1�{�4v���ӫ��Z�|� 8���絻�mC��|}f����g/D7{��H��۟O^^��E|Oemym��D�A&�A�oy}-N]�?͛OZ��jZ�n޺EF�!�|�9�X_�~Z]���MzEq�}~ƭr�Lb���㇯����=��H��UI�a�8�S��p�E��e5�g,YǮ�Ȧu� ���~�?��{'d�f]�ik�%����Y	��W���ZՉ(�{��0OCYD��8 �y��Y��9n]��L�
3��+�6�)���	a�m����>y>^`��qKͳ�q���`��䐩���<��Dh���;��n�e�ن�òY}7Eo��e�Y��VG�|=b<��:��g �0t�"��E��E��F�X�8�f�~�d/FN��4au��.ax���}�+W1�vO�@ȵ����q�h�4��;�o��锪H�0�2%ɒ��$4�	�y�fG\:7�U�����r6����t�i���w�*~�H	�V�/r ��w�p������P�d�ݾ���p������r�O��dפ��uӖߊ�O�������5e��fB�p��	���"�m"�F�y��*�/m<��fI*0"�Ts�寑��B�`�1�P�KXy�}���P�0�O#E0�/�ˡ.��g� �q�P�'�9�+����/��侱q��5�.���%
�1�� cQ�^�����+m�����!!Bh���Vl��6ǁ�,w�����Ŭ�,�m�nc�-0i�3|bZ.��n�&^S�'=������2*�bF�ҙ�S��X'�Y��[�,��h�f�cf����Yz�%��ys[�W��B2�6�0*��-�_<�8e�̢!D�M� Mq�H�i&�d�Z���]�pF�O�E�
�:��EN�����%ͩ^�Q� ���N��;};�U�D@�2���9�;�8%ɼ>i�.����*v��X+l�r�-7^n���1�V��֯d%J�59��WN�j$N	��+%R��oz�%6b�_�O����o(��L��^oKB��[������&@�o��T�֒P��%���B0���d|w
��
�Sl��$�������};t�f�jS֨b?�A�c�ڲJvV�D?�F	Ȕ�<H��m��&=�]~�v�ݽ ?�Ǵ������Ȇu��<ƺLB;��>�Q��I�S࿸rҩ��e2�=��B�0![#�͘/���WY1���r�C�[iD�$��Q?�B�ڹ�j�P>d�Џm���B�O+y�w%�.���K��馮��$s�G	�l�{��� g׾�V�^�i��d/5g��|T�w~�b��W7S�� ��	7���c�}�2����/�X�G系t��1;x'7�
r=�N���U}�����G��l��#��uC#7r��㱳�U�6:��s��|�2��ou넺 |��[��-W-�)�&�\�N	~ba�/"V(T�jQ)r_�*�s�T�QXE�J�v�DdJ�E9oy&��)�� �����l��H!1#M�P��tr>Њ�295�T2���ϯ��r\�����(���u�o���ټRhrT�Ќ������ �YF���"5L�ɵi�1�uH2tB���aL4��5����tk
'�q��w n�%���?��}�t��˶y��8I�H���_��ۼcip���~d�li�M�����'' �CD#)%{��
��>*?O�	H0��v;�Te1L"È�.ek�P�y��_j�Pv�`]ϒ���WM1�?\	�ufgb �`J臇d��q���vqP�K�P�hOF综�!}�K�(�m,�M��k�Mgڨ|��m�(i���Ϸ����R_����j����	޾�,�^J}�������5���U�:�+�M�k��A�5��~����@j6rß�L$�16�o��E˾���k�	Q]���E3l��닐�N�Sm�O���U?Y=1�-��Kt�V��c�4KX}�护��J1��sPg7�j����n�g�1?��N<����ֶiM��}0&1�q�6(~Jd����ط����9��)��8Ó�g8n\�N�#3�nqa��[K�V��vXhA��%��FK'u�ej_�
گ"k��+@�-ق]0��;�.��*NLB���SR�T#�WÃ<8�n���/��_�5]t���;�4
9�r���<�fV�#�����aH���ǔv��i�}ָ��0nM��U^�rVf�"DT��ĂqpV�_z��^��%���ʕ���ɽ;��	'��1ϗ�6@��F����ń>���GnѤ�p�!:\�d7��rT�/���ҤϨֵ�z��ࢄ#�دԓa�j�[�yfgW�xV�|N7��� ���h�a�a�$4)i<����}gj>��Z�&�՜Se?A�h!}X}�=�0��Y��(,.V%ǒ��R�[^�՛7p��%��r�������,���w�e?�ce�e��&�p��j�̰g�y�#vW�u"3�X�/r�pc�z}������Svsd c����U�ԫ����9_%Ϛ��|��RkQ�����( �72��Ez�|�_U���������F�M�}8��Ԍ��8�'���}mb�?4k���	hf��3ϣ���b�
uI���x�G���=��.�d����uAw�ȑ	n2��������O�r��0�oago��Z�u�*޼�K=�G�@���k�a1'}�'�<��E�w�z"`m�ˀp�V��Dq�ʝK��3��b*Y��)����,~*�o �O���In�f9�e��#䈓zݚ�~fw2E��x<��������g��_ݯ�F���U/+�RQ~S��hB�F2�W�K�#r�������S <�Ub�$d���l�Ve;��a��+���M��l�;�｡O�8�����������������ϧ;7�He��=gdv������C[�DDv1k_P��
d`�W0�����$8<,H���i��[{��b�M�k��j��4c�u��2�ך�̐7��?^Hª��<�w�,���Cf׏����(�m�\Č튂L~����\L�W��X�@G��hx�[|3(Y_����z�ȌNd�*��ܐ��.S�4R�8�q�}��ܸ���3�,w�T��?����� %g�%6����X/�v����%&7����K�g|��EN9D�H��i���9
�N����~+��
�0��J�Ӟ+�+���.i���NG§SQu#ē���2ua[Ȳ��yʐa%\���xiI`�1~P4:���̓J�F��Ϛׅ�٫M�m�n:��/N>�>ўJ�?a�t�؆�Ψ(@}�	�a�i���}d��;�U��O<�V���9W��䶊��LJ�i�1je��˓G��QE�ޱ"c|w��W����b���>"]h=��q�\��j����?�5k�Y�=>�ɶܳ8�����S��e����w�2����X�S*2��_��+4E_���w �p�\�t*��GP�V`<�и�$D
�p�i/�&��a$��BP�K���W۳U��ޓ䈚Q[��9�߮�L���f���rB�ēq��<��8[�MG����@�!r�W���pV}dn����D�yS���s�T,�d���N�§ᨀ>�O���ra�|����11�e��=��k��*˱�{2�`qC�vgP�� ��sw���X�ɾe�B
�nX���b��nv�¬}����[1K����>g�[Q�쇯y�z%�#��.�?bb���P��C��E~���br��cE��di��*ٛ�Ќ�i Z=7WY��]Ɲ��j�0��5 M�Jq�t.)%�H�;O��y9>Vh	5[v�U3J�b!\Mމ8k/6��ء[1��%�B��ֶ|x��8�\_�T���mx�����|Cv�D�c.\Y�H�^īkW�2��T�sI�tr�O&Ja2ή���7���鏉��y��$/׌��{�s�}\�W��-p�	��v?W�W���Ͱ_�j0�+5{X;��X�UG��� ��-p"%B%]����-̋w|�2�`��<j�pF�+�֕s_����Ņ ���ľ�D?�؀X����y�2�*w4y��`S���!�fߨ��bb��	�Թ��݁j&��yj�2TZ�s>�E%̨��Փn-ċa����*�B�=��=��P\�1�orP�è�m!�9A�	ΰY .���㯉�X�*:�̛�����Q�DE����/�[��-�WȓW�$��c)@ �a�T�Rp+�CLˎa�O0o^\T)#����CF��X���+E5G�����SS�I&*���Cw��;W #�i¥��6!\0ܹZ�N���$���Ơ��*�|�3���5�R�r��t�@(���}��ɠ?������}Bش��FE *N��m�5ZF���Ci�6�*���� �M�P�O6�-W%W2�"fb�\u�| ��;w�u��g�2�]��Y�
P�T�Ҙ�֒����n��jb넴[~�ޞ�x<J7�T{�RHq7
C�y<D<���"������ç�N�����أl�D��QLB����%ꂪ���n�0�6�j��_l*ԇ0�*��e��I=����M,V�:����U�\8Q��kL��_�����F^��{����7�L�p��b�q�$o_E�"���y�Z��E��x�yb#7_��mn�W�]�����9���b��~���,п=�L]2ޱ�����%��',���J�V�F�r�%1L5|C��g�,�v��o��G��bCjfJ�x��}n�tkH�Z�p��u<e"�#�E_SɭA�ܓ։�N)���,pz�;�h���]�(�?������0�����B�te�
1���s�豓��"�*�z@֖|UTҵL�0_��)���əqI#��_P�S��N[��ҩ�fG���|9�^M�����P2g��V�e�tw�dn�I�2��M��9��/Sw��G<�>�X�"|��7���wVleW��cx�*f���r¶yf��$��=���;5��:�4����A������_��%2/Y�I!/k���g/4���?i9�8���jSA��<��NxAU�����\v���o|)�j���`/^��e�k���_�;|;ґ�h�0ߪ
���z��^�y~��� �J0xqQ�W�380���B��@��<R�2�8N���2R
5 0��uab��zz�5S�8Z�I5P����CnUǈ`��b�]<��@~�Z�ŷ[z��p�N���˾�$�O�E�/��|�?���I��ɹ�P�7�A^Mp��y��9��d�P6��4�9���.��įx���ǻ]C�Q�q[{��!���IR��)�P��K�x~�%�oę[,c�����T3hWa}�;����#�Igڹl|���H�ߏ�ɵ�
y���Ќх{�ฌ��F��kB+3l���>�#J��~��<�j�8BhA6<mKHˣr����S��	��Ҭ[�s�p�HB��iN�@�3~ь^h���k�+�l�[ڡ?y�q��EK%��_a�a@	�`C)�}4�P�W@sP6�@���.����0!�4�ui�@�r��m�j?���>oaaЭ���
P�K��H�]�*����$Nb<��ל;���S)fM;�l�YDCʢEޚ�F�y��T3{O�|5
���]�x�Y���e�奇t��;#q0yO4W� �t�ldkO@����+g�����ch���xa���� ���7;J�sl�x���_�m�
�Ҭ�d�:��)7�a\bO��F�2�w�:yX��H���r�������$�U�u��Do���d���ñؽ�z�F��64���6^G%U��6I��0�~���t$~��#m�݌�*�3�0ް�B!G���~��z���%.`5n9S����lQ[Z�F.�{��^�{#G�/t�c��҃o@���|-�ݚ��l" ��O�5L� ���0�QS�HQ�I�p��Ϫ�خ�Fp!�D!ZNŰ����{cR�=�]cvv�w�n{��);>��<V�3f��
h��w�}��s;�;��6&�2�\�J^Q�Avr�\m�y��{�N��g[?l��ʎ�x�:�7�_���ۥ�Ќq�k��K�Ϯ�?|���ɷ`��#l��ù��"��n[�T��'�`xy�r���,������W���ssv?:g��E�A+���I��������Z������r�Xw��f�1.I�؄Hμ�u����p4Ai!Yi!�1��]���Z��������u�������9� ���1s�ʿ��-rv��S���*껅����%�3ܺf����d������w�n��ùӥ�6v����иפ��v(+WJ���8�-x��B�6�RG�X���Ќ=4&Ո�pv�]�򗻊����R0���.U��01s�XG�������py��/A �t�.�k0=���5MI:H��0�~i�Њ���y��x/n6�ܰ\���W/˝aͿ��x�g��Wz���% ����z�)�@�ӿmg5�j$�٦� W����G�Pʚ<�P���.˲:nq7AX5c�,��ks�	32J��m�Dp|���[reEo|~�h����Ѹ��C��0��{@r�3�us�ސ"�6���G��R�k��C�ΰ�'>�j῏���6��Mx�v����ȟ!�1��@K����RHЦN��]�/7ļЅ�k�2�bgWU^���ԡ�o�+��t|�0�!���[@U��d��I�X�[�s���A�7ee��݈�9�gOU<��;����Ƃ����c��[��2��x-���K�J�zt���e���m dF�8v�O�TR6�đ:��;�1�ϔU/7�B�o�9X0�E������n��lL��B�(-{2�c���%��@�W��10Ψ���^kvy�q�E�.|���ؤoRh�Y�e)ww1Ŕ�˜�S�J�f�kRY�@^��)�MSZ����H�+���$����:*���d1�R�Do��q,��kE�����@I�o��D:����!: w4У�� �E3G�ۮ�1�.e��Kh��`���a��S��\�4�8T��;��<����<����>��T��ާI3X��Q{Q�xT�#}#��\�!��w�C��/y���Y�E�u�U~ä����n�6��ֹW{==�c��pBQ0���1xo�+g����P��L�����}�+�^�.��taey}�;����-�7^�{ߌ$�Vi`0�z�ˇ���[H�m�7�>�I�D�I��ҷ��%r�6-�w+����!f
��2���1<+������e�Y��� �][����K�Wjb�� �Z�Z6x�9����/����2��K��6mM����Fș{<E��̂���K����vЩª��B�.T���TU�m�o����@�s��t9{l�EJH}�݇���n�&f#PP^��F�����ݓ���m~ ױ�@X-?�8u�<j:h�7ӡ���=#1!ִ������r���ϰ �[�ʩ���L��e��KP�E��:����uvЫtb��q���:��'�hYL�!-�X�({Z� /��y8S)�����8jVwB١v/��j5����b�(��tD~	��e\�z����B����jYF����j9����<����#�!%d�İ���+�r�:V���ހlf3
F̥�j����� #��@{�9����lj�fŒRf9�Z����q�!��!��6!]�wb@�vA��4��Q�@�G�!��z�@�g�P(��gK�v"�<V�������˅�̍���R7_��X�;>��L�D�
*�S������.	p9o�+V5��{�&Y�@�|�.��V�`-��#����B��0x��AH0w[I���?��%/,t߫��>�o��Jf���,�Y��	��!�gH�d1{@%j ~�'� ��N=J��,��]}���Q�hzupo��mGJ�֚6.���e!J�&5YS�����4�,c�tSK�Z��^m��%Ԍ:�-c&���|���N	�S�O�~���Wv�^�(R���y�3���l`���y.wNy��ϥ��*��s�G��I+��>2��ܝ���},�?���_oX_P�Sq��(/���	���J;�i22�h.���FMR�]&���*U�T�T�J�퀴-W��W�����e|m�̤7t���mE6(�SRd+lb�3NRk�\E�j/V`4}���yulp�|���WA�mK�;k)�����"&� �l��,�f�t����� ^�s�PDp�D	��T`hM�&mp���n�F��#����!s�j%%�����Eڪ1��%���ֆT#����Ȇ>�X.�S,6�lI�q<�o�2Xz�(���
�g�`���<�
��/5�[y�B�8o9c�w�˝�\�\"�;�Kr�-�ՙ+5d�ac���{�U`���jþ)g��x���J�&�<Pe��8�Uցݿ�?�G���,�/��^��J�O��n:�/r�]jd!��_���9��
�H���W[�!+��E�/�g:΄������C��m?���ؗ�ˌ�l�W�6�j�q5|�����Zu���P�هe&�j���dk�K�O9f�W�������!KX�J��4��{9&w~�,��*����H�[Xz�����)��@ޗ��-��65E���L�ӛi8c�iA�~@�����;jl��|f%_t	�+8�����w��s�WF ��kw0�.�Y�߻1!�m6��7fS�Ў"�>����:E�[\���|��-ēf�f6R�R}���ͷ�F�QE��A|�Y"w��O-pN>�gHm�;��40��x�Ӆ�G6'���	٭�c���6G�fv#ͮ,�_�Ϻ�M���0����/� h�ΙJU7�,���Ak�������<�Ut!u�P5�v|M���w�hϽ�ߓ�E�܀ ���{�>����'�]��G;鬲�]_)*�E\;�5��9|@�=sѰ�m<�ou���;�j��#���Z�>�]��2��`:z�ײ�W�����:�d��T�n 8�EE^F��^�j��� ' �p���|�3����>z���?�g�{vr��g�����}$Zη�N��~��oy�}�-{��QC�_�;Ě�Bhso	�Kz򊘦������]2`Z�g��Ϊ�:����ɐ断,��;���yoDZN�h��>�X��ԐHYz)�zBҸ�0��m1�.Tŵ�O}D�dK�������^4��NC��X�1��[4��ˀ�y��m�憌޺xG�?���*�l�?PCC& �i�Q�c��栙Z����*��V�x��%T^�hs���b��پ������,�׀*ѵ���|5 z�� Mz���d�u�Q�,�r��b�ю�
�����i2ސ~n��d�F��_��Fq�=4�U%�xAUf&�#�'��TV�[y[��ˋ_`宜!]�F�?گ�W��j��Id�&Ot��}��ꂈjM�<ŖGC[@����K �A@?v��r�bYh��Ddo�m�ktOet�m+W'j��$y��uSh[~���_���9����𰢱���U�^D�8�T�MbdJuY͍��eK@\\p�anN��x"�y�HJ�Q���5�SS���Z�?�ɗ��^y�<����29���!��Aࢋ�M��C�J�3��)"��>�8���*j��oI.�q�uβMs�3�F ��3��[OZ�5	5b�Wɾ12�
CC{ �a�bK�{a"yo3���/����?[��o�[���c<E�~��)�QΡ}��w��>2��@���0�+����s��e"
)������8N��FC�,,��]:~�l(Y|�����/|5Nf��Z��Î<��gR����z[e�k��0I�Ղ��X�بʇ�, +�q2��������R��kB9������Ϊ\b���Dʺh���E�A�Ke�{'אw�Y�Wߝ������׋��cs�����22uaZ���ں�З~	���v�5|�T#~�M�+���F�M��^����[[����A�f�����֝Ҙ�¹�G��֝���
���0ghxJbڏ"�n�u
�� g�eV��&>}a☛�k=(B��z���#}�r��p]�9����nm��d��A��q��V�<=B0���	mA�����b���T���XhŦ����P�Q��g���d;�e�+tm]M㠑'V�I��V�g�.R@$�˯	�$���V��,�/�d/,���p���ھͷ^-����=$��Ok���XH�H��O֓X0'Sm�֟|��O�Ξ�81�
�.�Ӟ>i(F-�V,Nn����?�c�"�byN(6���2�s`�v��:`�K���Fuӟe�m�A묚E�a��X@GJ�����B��e�E7,��t�T�Ƙ��>�?��d��W�l腫�����=�z�����yEt!�o�GJ���l 	2&~M��c� c0ѩsk9�E��J��M�o���U'ځ��П��J5	�c]C4������
�^�ϩ�����~���v�/�d�4qn�E��O�X�+~E�z	0�3ߋ1l<�7�LI"�:��S+ڟ�!��4��jӽR=Y|�Ӳ,��/�^�o���H�-k�~�y��a�����zZ6�?;��9��ůt��Yfy=���V]�;����>�`�<�U��;�{3�!��w�B�<wu؛�8W��~�����?dεSa(�p2N�4�x�d��������"�� ��Q[��T�}����gH�� �pu�c�aQ\��	τg_=����5�����	̍���h@"�3�F�3�Ը�L+yDrڇ����P��n��9}���EΫ$�(u�����j�{� ��E�}��?s�C_� b��@��7���J����O��R��1#sH>3��=��0�(���>�fq,��13�T �N������� #�'�CJ��&���.���0z��F~��}7ͼ��HE�ײ�Q��i�X`ܙF=�M�vw���B:?���W�P�ذOä�lx��<{�]x%I��H?����z�q�#I��q��U�ш{i�m����#�fC�Uh�W-��~YZ1��ף� �r�I�uDm�����5ts���MfH��ä��/�D�]�N��G��,��>t>&�GiF��D�i��2���p�5��t0ێ)���τn�;�&���#a���0��=a��Y�F�6���(���	��.Ҷ\�\���1��������dc���7諢ǣ����1"��8�̇��v0������!�T
L����-�Qj��o�4�r�F>1��(>���d��`�;��A���2�h9 �8/�s���ڐ�@�-�� ݚ��nj��m���_Q�[R �F'zʹd�U��L�hl4�]��3@(�xܬ���w[~6�/�f@�62B���-:Hi=�XhY���A���WH��>'%�`�Ow���H��ڹ;���yj��ޤ�6��V4ز�Bgo�r�GՉ��
ÀѴB���M��Y(y/{V�:��B������@�J7�-��� [~��G�������Q�i�>a�(�޿��sٙ�����
���A�qb��	�$%�]9�5��R�R�T8�,��	Zđ�����˙R��x�ӯ/��|樳�.we(�,~�<\�ٛ��/~d��$�uF,�I������2��w}gA���f[���Y5��;�|��A{���@�y��"?�^����S�*�	�� �'���L~�[��H�@M�WX���~��Y<7��N]'�Ҷd�	�w���jD�ޘ�)���j_��J�i�ٚ[Gkn4�z"��[X�@~@&�j��i�^~���줕�'��\FBc	�nƈGۂ�1C��N�[1�U�����^h�yf��1��R��e��$�r�+�����LQ�&ѹ��2}�/����*�f[�i"d�M��n�ŭ�d�*t�=��	ԋ�R�/�#��� z+�ӎ�D��ֱ��7	��m�0������� $'�d�=M4�b2��EB��۫����c�	�*�)�E��JE(pA,/�	a����WBb�6Y9��m_��K����U^6GK��u�����ӌ̡�t�#o��˙���SXu�l�WTM�ȭ������ݥ�.>ٹv�n[b?��t��n�xr�K��3������ʽ��K�t��3��ќ5y�Q~��J<�R�����&�#> �^*g�)�R_|v:�W��&1&���K��D�s$9e�}��Gd6�/��R%�cË.,��:!��	����z�������Z���66�b/�8����:�/��SqŻj4��5�`��
��J�@�D��(�(��x�	���m�\�fk��_��a��	��w<����G뼈IG�B��=>?`��̕/�	~~[������Ҕ��/�I�P�q�� �"��$�a�EW$l�s~gh���K��<���e�ئ^Y����[x/���eM;����V�΀8�寧�<w�G�Y$����1{nDL��n���r���b�r��<��kJ�����������6�2�)����*�yT$J^�/��?H8���lH����"��G�����Aѕi��w�����p��ٛ����/ZX�f&J�k�s�yH ���vdc�*�%_�t&�|u���v�Е��eK�tO���J��B�M�hHL:���6�ѡW$��CIF�:q(��]ٹpF�X����G��$˨̀��Fɔ���X�^�ڷ�O���w���|�cl_��u\���M�Zi+�0��9�5�����X�����o;e����`ϐW�w�X`!��8�N�֦.����[9�Vg5�/Sr�����U>=��p�+L��~ӗD�D��������q�ڛfYm�L��3��tBg]دF�N2Ç/o��Yt�'�K��6�+�~aۍA-	��#vQ��G#d"����k~��˳�+[#T>aa�^m̈́�Xh�v���������ѻ���h�Y���oGJ�o�>�8\<�����E���z���:}���y��J��b]]�7t�~j�uGd��j�f"�>����O���S�-���c���7!6W�/�M�M��.{.�Q�b��G���g��� �#��l�0�'o�l`�|Z>�Pz���|��s��T�6����#�u�i��t��9�4��m׌��c'� "z�c=�)�[hQ��M-S���Dӝ��go���5-K �Q�"#3(j���Ȇ��`�O��~bz�z!� ���T)�f�ӄ~��[x|���3�q�x��$а^_����N���o�J0^�V[�������}����8W''M5�g0�'�����1쏞)���I��q���<�w	�0P�SzY��2ޕ�([4�׸�^��n)vᓽ�Z�7�}p�ܶ�ïh�o��Ë�A������w�StfI	�Of�2W��G�j�E[cVsPG�����[J��3�{_�����R>s��ɋ:��eD���sg�)U���s�!˰�#ky����Y��<��~wۦ����y-�s4��s赤�_[�_M�~292>�7��0&��9��f�{�"�듳��L��[�p~n�����ǽ�x�[�W��)J�F�g��m��&�@���R����)�������6��^����ɷ$0{���"��- �/bk��lN����b��X�,�q�SZ{����]�Ǯ��WF�)I�u+�-q4�5ץo٧VF��s��Q���04����D���뇱X*�#9l���i�O���ܚ-<��Z��z4�����s�?ʀFb�8���//��3�,�g���
���.>Y�`�^ a�I��:C[�{��^#�h3O��ŧ�ج��O&�[z�<깾�]#=��l����u�/��[��X���!���!�}�>�)��)�8�Tc�b�����b�(�����A.d{$��|���JaDCf��Ë��3&9k}��\��t���f�}y,42"O&0yC��B�[F���&���K��[I�gYL��_����_�֙�W�9�6�^�s#���<����R7%QD��T���t��Pd�I�����f+�)R1D$;ٷ�dϖ쳐}��3f��<�������_�y�s^�9�y�\!B�v(�Ζ�6�vWK��ԁɞ�
�1�O�wMk\ׅ��4O�Z�/,_(�в��,VR��ϧ��^���O��~����B����#�� k���ɳ��XD>�=�?�rsJ{.)=a7�R���8�X���j�l QC����R)�R ��u�iT�����DXYRT���;�_��F�ޅ�;�������7���\j����U�r|�-�f�#�_w�h	<�f%mRa�+c��SJ�/�����I��}�`��/Q �^���b����J�T�" X֕`^�ew���)[s��:ߖ���/�ǃ�<�vrO����:�� �'����3^Z�1
�E�����mmǂV_6����\��j|���yU���PoC���:�)A�� ����V��)!����$>���5�yWfϾ�c�,>�x]�t��@O���3 �� !��\��2��7S�j�d�Y>��S�D_Es���	���=%u�G��Yo�:������M♜�֖s{���%=?��R��E ĉ]���'���s7�x2`����&Dc�����a�"�$A+�m�]��<Z�}�as�6[h6)\�+�NM'�����\�@ᦕ<��^�T����Pgq��H�Y���/�3me�9��ub����;t1RY�4�{7�����bE,��n/~���!���!�9�#�4�h�����V�#��!\ߡ�ǲ\�&0of:6+�Q���J	b6����U��v�i�������+�)UN�i�\1�vR(��O�.`[E�/�$���s���jȲS{u��ԿQ�Β1���n�CA����|z�O��Ȅ�r�Nq<�L������P� �ݺ��(��u�y%, ij(��g��H�}��0N�l;��3���b�2nh:+� ���W���f~y˅�}�kr;�d�
�� C�ꌸ��f��8�L�~��ވ#��5�zՎk|�9 �Y��4��G�	�-I��BÒ�J�ф�3PU��c����'�$f_�=�.zD�B��a'W^�������v��̔�d���3r��uG&��Bֳh�D8AŒv�7��b�B�Xc��Oh(� �q�zz�_�X�� ��O*80�~4�ҮV[���D2�n�#�gD�|q�< G������.�\>03�Ȩԉp�ǲ�s@'q��Q�3h�����G�6�=�Z*��ʚ8��B��&�4T�;�[�8�м��ͧ���ȱ�c3{�UX�O�m�x�R��/@��{�[4���S������;�摪��G)�/�$�5��J�l⏠T�k�&o���c74���V��罹��U��t
���ૻ��5�IT���d+�ѫ	=�jn]�U�e.�r�2�����%����i�O�����ms� l����?�7ڲ�X�'K�>��W�{)�Dv��)u3P���^�A��Dh �c�����?Z��;����}���r�@y��X�&?ي�
WE��7hrİx����%��S���n����i],0�4X�t��re�i嚫��ָD��ʕX{��95�*�H�Ɛ�h�dO{���^��5�ĳ�����;9Q?�W>��*Ί�l��2��IE�8y:�M��Q�jU��������I�y�<���zX\�b;)�]^�;��b:�|V�%h���@�g={z�}�/�C�c,�����g��Qaw�" e��5{��͛�I��S���B����HɛN%UK4�@�����AO/ru9f"2�ψ2�}g�
��h�n�<l��N<�>�K�I_2X2�J�F�T���@�W�:U�$9ܪ�M��4���y�����U2��	��H�}d[�A�蟾�͹2b�%�.�������!���!�=�P���P��2}>(�ZM�\4@�����}��k�Ϩ���&t�o[����SL�h�%��Q��W)	41���ݳD��%	[〉1�I&:+�O�	�{(��X�33<��`�I8�Yx���R���0
!��pQURĐ��f6%s�h��@R<��b�P���_����;<�1��|��o��^��z�w�F+B����~^�f�'�Qi�����(���o��Wt�"��N�
p�e�\��������u]�v����ɋ;�r��t�{�#��r
b���a<�.ݩƹ&��<LDl���3#�Q�����e�I@veʒb*ǁƏOF��Z�t=�ƥL�_GEs4�k��]H��Ǵ���9ݯ�1	)���}P��9�V�|�`�Pm��vS�#����@�N�!�yH��Oם��7��/� +���㶬|�}p��
�5�WF���mg�J��R6hIH�����8֓����yqu]`D쇚xgD�z�64.AE��,8����3P2�;IX�����;[��:�	̦�@��v?&�~>�vKxD�8����=aA��Cm�� �'����]-ڸE�q���"sA�Z���g��V�cv���O���s{��I?H���'��82�2��~o牍Ev��VwmҥA"�)ԣVJk���Q���g��c�ܐ�B������I��=S�C���@��c������q|��J���z��n��zG�'ڻi=�q{� !^�B�j����՝x�u��ߴϔLp?Q���r���d��;7��n����s����:	�1�	(2�'�E�O�?����7�:��uQG�y&Y@���]��F��+�ю��t'~��f6��SR �[� x���;��x�$[ڝ.��͙��!Y�(ǔؼ��;�,)@V`7�O|�]m�ub�'f�)������'ߙ����� ]�����U�X�����
k�M5�wz�xh8��v(�r�=�p3��W����`]�@��:���KxW�zu����q�@�2����Fj��}���GP�
i#ϴF}l�t�:d�{��� ��PR��/@��ˑC�I˄$w>��"�
��&���xu�������<T���6�~�l\j�����v���������7<�.5f�)��c���/�͸O5��	\y�V����4��5_E@h�W�G��=�ȯ��gc�AP׈��"?��Z2}ZΏ#��4e�td�С@�f3@˒���*в٤?L���?U���s[%���l��\)�˨M��g�&7��*)���t���o:J|����A�D���qj���`L���4&���J+/�9A���`�%�e'`e9*�i���։��NH�\�\�W"�iӬ+΁[@��[�iY}}
;����� ~>����W]z�4�p�2�؄��C�:�����=�W��Zn���,J�]��W�������Tt�v6�#$�.a���/��r:���jպ?"l>{/EL
�AK��\АR���%@��k� PC ?��`e�n�PE�.B;���>*i�G��7����P�@�6�j�A}��;\�xq�r�_*MW]v�j�ȟ�g	fF��?��|L����ߠ �.���5���V4�^��u$N�MM(I@>q(�x�d�P<Ю�ϛ�so�U�ۖM���l�qM_e	�g�XL��q�*H,���=��ϣ.���B���:T-���<�pj�*D x^�79�χ�ε��W7�k_Z��n�1$�pRjS$�� ��oau�w��P�|����n���*��ó�8����B�4��i1�{���o�B��}~�Wܥ���������**�6�	�o�a�9,�zZu8�:F�u:���>h����]�\��O�Yih�4RZ���S���S��,ޘ�/���>,|�6@��ɋ�c�p����=�x=�;@�����3�|�=3��랠V��{���������0
n�x�
��
�e�"[_�������%���ߢ*-l,��@u�������(�=�2�a����[��6vhxh�P��p�q��CRC�2��#7DN���E�QV��o�����x����l�C�W���"d���@�9�ㆁA3�2��4���y^��@tG��H��'���C��@#}6�T2jt�mh�МS�O!C��޷�,��ing[`k��Gj~/�	�[�$Xs�|��x)��c=�GB$*�hX��ѱ������lE�����q�@�b�wVs�^O����"P�}A�)��3��;Ra9���w��1ͷ�T=��A����n�j����\e���Es�
�ҽ>��6���?�0�p�?�6�>�j¸�r�H���S��j��rF���@`�77���V�l�-�+h�إWdj���6� ���a�%� �%�i1�$��nJ�',OO ۺv�� 6� ��#�_�{F���ފ��y`��fOA�ٔ���Cf����fx�,�Xu��)���v� ֍��z�x��̙�[��[��VwS�_"�i/$5PG����7�Ҋ�P����f@ӀŦ�C�P�����T�҇����Y��)%��-�˵���v��R.�O�a�ˆg�tj��DJ}H0Nk</NI9�a���'�h�6@�a��xQ���)�$^���
��:�?��[�!0�����\Qg4�CX�
���x���
��y
����p�o�$ӻ��0�ة��p{/3A��������.����--��w��u'Bu*��5Җ�m�� }��kio�]��ʺ~��0U/r��(2\pPzA|������){������<��d/!S�tС�Cm���$
���ܣ���!v��f�#Ûo����M�����e�4�\{ �A�)�����}�P���T! �9��J���OEG�ʭv�;ϳ��k'5�9�1�+�D�a��C���&�	4j$|b\IK�8���y�Ԅ���)t׭��!R�7t�c��O51o�l ����3߻�P����G�42|�ye3��@�1ʽb���(vK5	m~[Oc�"٨���[#��D*J �"�h$��Q��l� �U
��Khxp�'��4��T�{�v�o�X@��Z1�F5��l{���	�g�3a���k��C>��5�Ng���&��i����ģ����+�@�GH�Ym��jt�$��*u'��t�> ��h��m^|JשCٽ n�*#G�\_X���ɝ�(�8O�Q���`�Q�X�a���|�-q:�ku(��������~���/,��=j����Q��Ts�L�aef��d�;Xל�g��yE��+�SE�sV���do`=#u[l{��r�~6?�u��`�8L�>}M;��7��_�Q��y51�?qX���*��A�B����!�S܁�v!�jx�h�m�2�;�l��x ^ �6| 9����x6�p�����@�R�٢�w�:Ō{�pK���4�ԂO����R��ii?o�;�L��CxO���o(��S��H��&AǱg�3�w��eMI�O	�k��$���O�I#���f�	�s3�NU���3a�"
�sr�qU�oKܴZ4s����_��6��n�c!����������4�V�}�k�F	6Rq��Q�8���J����~��O6��� �~EF螸��>�D��+�吐AeTq0��FX��
5g>֞b��i�f�ii�5�II�E����.����9]��&�0�;���(�G�oB.���C��\�+z��w�tL�G雧%?w��}�7�E�n��Z�fc�������CQ<b�Źs��5�;Q���)���-��J68�O�]�f�E.�U�ᛣa�a�}����R��\��I��YS�U��߆��ޔ�U �䴒2�\���VٟQ���
����Bl&��Il�w�݅
���JI����}O�O�jQ��G�%������=g��~�JpRA�L�i3�N�M,U�Q��/�\�ov�t�hfS�C,�����[%�TnUE���p�u�m�O.��s�]Y^�ڼZg�)����V�>I�]�7G4�F��P�����A��oÆ�p�����C;�.���T��x�|I��ν6p4pA` �>8`�m����!�.�,ՊE��9<�� �Q�M ��\�I�W�q�$}��;n/��	�"�|�e��2c/�CYo�����uN�,TO[�^\�S�\�}E
�u\%���^�.ª�M껨�Φ_.�*jF�P��/� ���C����$W�N����YH���>�\Kc��a�V;5���\�5��0�����X����������chj��E�6�N܋ E���Wp<��%�K8�3]��OKr�M�g��T�����"FK�w���Iqmsu���n�8�\Qš�-<b7ƃ`�K`�̙����Z�Z=�����U��u�F� Θ�#b}�KLY��±�/J�nH�և��}��[&�w�+G:q�%-j��B�	.�1_����6U��s�}X��ϟ��ș�Z�������sm��#�J��iH�֖2�4�<ɫ��ˋT��ZG�PӆO�����A�t�:����� R��s�}�(�z��<ϗ� �y���%��@�7=��6$&�B�^C�2���������mJ��yLb�DQ��|���5r�?5��VT��}ec�)��,
�S��Q3?W?���͘��Ӕ�Ǌ�Fj�𲡋��l�����)r���b������5M��o����z��7H��ٝ:�AB�C���a���g��O��N��~����pY--��~K��G V�<4�j���7g�F�eZ�,z�� .��:\\�g����P���X�Gi�1^ЍƗW�L�������:P��]��!���2�����ȡ�<��=o�������5G��ҁ� �
y{�~��ҿ@讥����#,q��Q���4_T�!j�G:f[�/{�)��v�}Dc��1
G�����w�_�;����j
VB�5��HT�Q��1����^,-t4}���=�^�i'Xly[���ף�S�:��^P��������i��Tv g#ⅢNq��N�x�{n�!�d�;��?�c_��3��(�Vޅ�}ӊ�]I� }��M����`�+��2F1U�#Ԓ��5]M���~iE�K�p�J��<y1&<<q���!����O*\~n<3��~n-�m�3�,k�@�e���8��%�B�n���8��p���an�V��d�pš��c����q6q�4��	}��,殺�-�)�/�� ������߅�מ�M]��n7���W �i�4�:��RB�q�lK�·�Sb�}*�n]�Ib��0T輁a=[L9����h��fF�o��5���۾$L�=���S��<g��ؿ|W
1��΀3�%0�F�������G��V6:R]�w��\r��޿$����_���
3�A?&��EQ5�����>օt��ofF(�;؊�JԞ׊�sS[y�/���ˡ[�x`�~j�7T8xB�\���C��잜�0w�t�`��p7�]��*��O���&��O�u0�\7������PY��B�r>푁Q{}c7wA�.�4��!�������y����j+�h�۟x�s��|t�;+9pxc�,��T���� ���\�m�	��G8~'@2f���F�A^���4}�{���m�X�L\)��l�S�k־|
b~{;���/�c]8i�4���-�/�<�9��W���~A\X��ߎ�}��������6}�uzz��I>
em�L|�w'7P��;U�EV�-|�m��?`��A%��v����I�?H\`h��o�{�ݔ�V������{��|9�2���_�l�ՌT/g�-��6�o0@njC������F�`��No�kSU �������P�,���l�%jG,��[+����RkĒ,ga���!�������1���z�Kd�� �i��#�vS��P(������}N����Z |!�E��\���SI�k��|���?�)>H�4�"q�>/\����(��9(rthw�p��%Ay��y�W���ny?��&p(������+�׍�1�Ν�!Uf���g<R�h��	v����<"&M���?31�{��~I;�}�ѡ⧨��Kr�6I�0��q/����2�d�[]1YY��3�؁]ZDP�d~�6Ū�hN)K'�a[����
����V	��3n�JouTo�$::����N����5L'r��-�`�ڝsm:@ld��h�{I�"vJ?Z���m�DT�.,?
���_���/`�씦���o���, f�gg�y7���SF�j���*�l�r�66Phyf��5���<���@ø%�h�u~p���z�f�4P��?�c7X�e�|��CVw��G��O���+�y�?WȾޔ�]]��f��� ���F
0�1���z�:-j�����S�~�U�҆��/劃{� ֖X[�Lc�<�jb�s��FH��̿�/5�?��( Z��p��4���-���L�o��� ��"�?-Q�(y�����{�NXcunc��8������b�t��D
BHY'�PJ����߫9!k �m�Ԝs�%�q_�Wm*\�o�i'���7���
1��Loi��-M�����Z�t�Ȯ�2%t�J_ �%kذ���΋���G�.7��S�FV�\�`��׺�R��qM	�zI�қ���~�Mu\��~K&)Z�m�,-ψB�Ґ��R��_s�%���v���_�c�wX���q�i|J�r3�~f����D�r����l3	<�}�]u]MZV��h�����?�>#2��n)���$����5���į�{ye8�:/̳�3���t��ܻ�(�.T4�>2,�$�6�ͬ�w�#ߔ4��Υ���z���d������>�]��_s�3��� ��(Y}kJb�]�ߪ��N���L8���U�d�K��q^+�C7v�=\����^+l�X(n:�Ͷfw���+C3��\���]���߸,`������,Ҋ�!��WQ��B���G��c��=���Ш���ŷO.'/c�J7��Ԭ�������j��ԭ��R5m7A�>�@��M9����цjk]���N���W*aP��% S� �Nx ;�G�gw>�>����y�p{[�!���!��ပ�WOz,�(�T;
���vv���dI�V&"q9�86Um�թ�9�ϣ�O��y��j�R�w�A����_�w`�a��:���g�� �s�nx6����9���jF��l`�_)��
���\>�ߠݯzu���+
���=��j=��8jg@�Z�ۀ1��;����f=xD�CV�G��R}�1��oK����A^�ܷݔ������5f�f�~n(�`�kT�3ս�4l���vR�sX��/�i����<����Ԁ{����	6/�o�����2���,�țwhM�?��<�,�}��=�*�B�Nds����È��5� ?�N�l��ǑO���)l@1���/@�>/�E5��+�Q�ʬP]XO^��?�#�V�d���Ke��:�,@`�0b~Iخ7�[UrA{d~/Z�㋟��s�	�%��
�0� ���S���x;�����_��$���{&���r�|������z@�����^ؔ�{T�Ko���ʦ7�`�{{�}ox��ϡ��=�0�|���2�z��9�;q�_C��.��HZ�RU�X�v�IgU�؉_��	��i��������+=�?���Ud/΁G<�F�6��FJ�-��WR����?\�<�:A׷���6{�I��h��nOߺ�y�9�N�k��uv0����-C��^�2NXy���P�ls~�r���Oxx3���^p�����cl�d��<ĬeH|�V��0���=��	yX���!v�p*[]<��u(�=�����u�'p��%�o�Xko�q~N4����oI�)�u��>o�����w��7/$毓j����!5-�+hP9�8���<�� 	�<����@�Ojy!��գ�Z�Fվ�ZZ{��0��]��YH�L4�K�+����)k�o9��Ԛ�h�;b	Ɏ9X��;8/4~5�����i����&�`9C��������YW>ffda�M���V�7I�`1�H	�x��	c��� �!����	��?g�֮.��h����h�,��z��{&�͌/8	�y:]�3W�`��GwR��)gؼ��:�b���GdG6�$��1u��jR�7�-�X� �rk�iŀo�kt Ӳ@��OS�-~Ҥ����rZ�2�]w�f^@�E�!�^q@@>��}.�It����ԝPT������@�M��/K�V�2J��s݇=�cN|�́t�7]�U��n���:��إ�}�rn����0�qm����=@�i���z�QV�� ,�i���R��r�d"�8J�*�x�.sDR�hŤ�a��;8x\�'���8��>wWm�Dy�R�&��|c?!�,�Mn������E�ض�`����b�-L�
uq�z����g��)a3���UZ�=(x�g-���u�x�)n��D�I2���}�4�[������y�?�ȋC�>\
C��g8����,W
>�t� ݩϬ���~2@�<�&vX�Tf�^��N�`�@�d�
$[�����s�X� ��;v�=�s^�#�+$��G��\�U@M[�B��1��� ƅL���&�%ʐ�g���d��c�o��P�2;k��'8�G�+���]��T��)��n9��ڐ����[3Q��,����0l*\Adb����h���5��[N��|��SC!�8���V�/��Xx�����'ކ��/�U�2'���2����~��AeL�R���/��}վ2�����@!��z�૩���9P.��j�#���*��������j��lۍ'�Ȟ^���ʃ������d5ۅ�/��̦mg�+:��~�y�S|��=*.�FM묖����,��!��������M�Z�唭�ޱ��g�J�~eۅ��̥x`R�J̡����:%��s��1w��؅p�e�}[����p��{���@MM���D_cM����#�$�M%��ʲo�m�L�uA0p��m������c|7��<�\���r򞩮]�b��$6��ۢ
�����ZuSqzr�Y��	�A��W{K ����լ���sx�1 z�ǫ�������I!��7�/0�*�ت��mguϻ8[}K�L����O
�<ɟ��I�n�aU.�s�$����m�z���ک�����:�q_J��̗��8�����<�?l��g�a6��Wj	��7�'���z�謵�V܅��>�;��n�Ĕ�����{e�$��c�K'((�ɢ������m�*�և�c�2G8�}:���H2-�H���.nj����ܙ��Ofo�]Z�b {�[Jr͓sjK��"��׮�O|#bE����e���]���]�=���B�	�0��$�J����Y�����̙�j�c�X�aN��yX�=�A�p0��z:O&�mr�z�]��kewi����-z�Y�=绹1g\l�v1��*U�J*��d~r��\�����]��|J�Ne%�k3-�T����t?�և��-�˙�1m�u(4.�C���f!IQ�4�N���~;H���no�0�/f�l�t�n*d!W���OR��eYq15�~~]��V{��y�,�Wȷ����6��w���=|h���V��B��Q�D��[�c���$m�*(���i���5tG��ť'퇻���b�\�:ۥ��$�$���>���]l�R� C���P�#;zf�`j�@�K�J����$v(P�Ӥ�ec��M�X�,�}X�)@���V��*�����}���<���I�K�QUxj���=b1 �R܇>RO�������	~$�"�=o�CT���F����� �����}�������n� �U�� ����4P��<�H�C��|J�E��z��;��dq�Q'�P>�a�q����&b���ߺ��m�>� �T��r�YZ7�_��c���ɀesaiKX*�Z�2�W��\<X�K�|�[5��hA�kHp�4Λ[�ٙ\����K�~4>w�Uv�^��0�Գ'�X��c�p��GA��H5���G��ځ&�h�s^�\�G�1m!� Q��j�u�%u�f���yi��H�EV�~h�q�8X����X�؈�fpH��u-�|5��+���nP(T�T[y�cxqG����ωS�^-W4FJpc7�9�1�����xu��Ǌҙ6��G�p�T�a���9X�W{���$����vo�zs�zx����)P a�έAC���+�@b��F�i����y��w 2��K��z�D� =WE@l���#���4pe���
�P$% �F ����;��p�e��ʓ6��;V"{;1W0����$&Fzk��Ĭ���o<���e�`�򱂑�:��&�p}[/��Sbsn�4�u̐���EFH5Q"T�N؅���3�?�Qcl���A'Xt��H��$kV��"U�G����W���ݼ{v`�R8(lŭ3��%c$��eH�P��x�`{��λ|�H3MJ�=�~�.\t����R�e4�4��e
1T=�����i�B�[�E���e:�1��H�ȟ����Lq�upR�-!�<x޻��x�����U�w�<`Y�����!5�vCx+.�I�_�����̈� � ~ǭ��ndg��^EV8�͘V�T�~���)<Pq��p1���c�|qO��A�?�A����[�ŭ��T��Y���I���K5ȴ7�_��C'6��^ޘj	�Ul��[S�T0&h�=�U���0?��,[�6�/��H����1��/N%��s+�~Ni�W������X��7�U���Ej~oZ�P��Ф��,��b#�(�q� �s���ã+32��>��قe�Q�į{����w�ݑ�o��#'Z.��~��Jh�R��̓:yӫ_�4u�ټHÕ�e�MU�'ͼMR�Ԓ�0�rGT֧ߺ���1�K�-�R�ܼP����.�F�ĭEZԱ�[�ל����q�W���}�OY�Y�H�6�I.�>���#}_+!��^�W��E�qq����L>V��_<"��J���?w������+�x��i}�sP�i<�'ȟ����������.9���iC�>"��[�ދZ��X\�+���?���0:�#@I��;�f�X�Ԯ�a�r&Nkɷ��F�D{Ֆ�na�ar�WP�X,�JT�顰�Y�) ;�8�crz�H�J������y������XHQ������20�1&�3��v��H�Ģ���O��@ 䧀Tqة}+�բ�3ϖ�ze� Ӗ*i�/��e���c/I�)Vg�&��L���Rvj"�� 0�Ƚ =Ǚh�����V��jP�QWY�	3��Ϛ]Z�g�����;ws^B�)J�gʕ�v�К�{���u�',h=Gm�״bG�RY2�+�]p�3eGg�J����}|��7m���gGͧ���ڝK�ؙ�o�%�
���fI 3��9�P�p�� 5�9a�T�����%�߭�~����y��Ì
j�e����zo������xN��tU�!���	z�B"���z�䴖��DX��>=�I�����s��02����ٿƁ:�����#da�ջ��S׻	o�,_!���j}z4)i 4�<��>Rei��2	F9���L����)m3&�=��vsP=9�]���d�\�6pO�L�g*aݿ�J�&�J?����D�x��Z��d��Y�b#q��
�L�������54��uv�^jSjb5�)!�*8u����de�M��L�痊NQ��8�T��J0*>t�����;y����Y�RF��&&���������{S3C�7	��N�}Փ Cl����!�w������D��⭣s����w?�vŨ�p����_����=ѯqEANh��p�˘I�`Ԃt����Q�{�};���A/��5�eTBc�Ă�qk;T#'T+��ƶ����m��9١Jz��r�$�#��ܵ�ǎ��׸�?E���q^�j���,q���Y�?��c������@�P��i�vTݯ����]"�����R{���Hɒ0�y|2s���y3�TЩ����9�g�2�s�.1�?U!���o� �)S��9�GD��`Ǧ��Rgu�wl��ρ��-(�mw�����)��DP~J����h�c�3�U�L�{Փ�nhTK�q�K,��2˫Q��������c� p�[BŌ�o�D����%3Gʼ��Y˷�Fo�K� H�ޭ{�#4���D�vz���ըa���|ٜ��(�����JbC`ay��rL��(GB�>H�c�� �SV��U�R�
���ß'�Y<{����΀O���6&׻��Ӆ�Qbnb��w���,Nƅ98G����5��T� _?Y�9�qM��oٰ��R0W��VW7� H���RA�����o�S�~�Ο����g��x�^KY�����N��0�~h/����0¼�ْw���=����|uD�>�Ⴖ2T�&pQ�HJ�dt�T���)<e��b1V��u_8� A%�R�V�?��,~�v�#�pe<���Oʺ���/{�}}1�9���u��ֶbBf���3Y���bK#g�"�s�k4��o^�A� ���&�>:�=�	��U&X�����5c*�Veb�`	�Hڼ�K�n��@��|D��+�똑���������Zyy�t,�*U��p%���p?X�"?�(�?`M�A�~h�#���E�?X��LJ�MI��Jг|���JeA���Fb��|����6*�DNefż ^Y[ՁGc
��`��KV���,91�E0@0�]Æ�R�MU�H�|@��Eo��$��~g��}sp3�XY���kE��t�%o��	x4=�Z\�h����@���S�XK��^5���2j*Ɍ����С��_����B��!��J��D�n���@u!���Nּ9z|>���&M�u����0-}�����z���p�&��Z�P����*Լog��s��e6�\�����H]�CX�~�.��L����ȼ�g�n2�ﻖ�Qnh�Ժt&�.�qh5@ �_���Q4�����3Q�O��1�
����p#f㏹��\4��Tc%�0F�>�%�\�)YI��q�^[L��5�EG��֎���C�w�(��;Kl�����ɖ鷛�qo"����v
J�C���F.y?QB�X�^؎��:ή[`h����<4x�P�Φ�<&&�yI�[S��/aJo��OiE�QTb�L\V��{rG��|�����9�� �	4����vCW�J��,1�}�JUp{q�7�M�%�u��Ҏj��L���=�B��(���z9�y��{C�9�j)D�=��/m�F�G���/�;�x<����&���Į�I���lbQ�0�r�*Wŝ��<�\0��VX��Q��g9Ce�-
ì
m����T˄���FC����EZY@�����;+/�y(��N��&�&3d�8?�2�ȅ*�_��%�'N�	B4�|)� Ii��
;j��,��̨��}:�08��ܙޟ�7�G)��`jMll��'�[;��C�S&3U�;��n\��2�G�8+<����b>���4�j{�	�"�݊��37oٖ'j�C���^o�)���nb�Q���2(�����U6�W��e��i��89qF��I�5�E���.��P/=�P��Ul�x�J��t���hD�X�EN���>�ș���\�WXۇk�~:�{Zc����tC9c������K��5���N�C� �(:P8A���(�R~��	6��Oy!-�3�(����9#dB�F�D�v�s�`��A�Ml��VX�'~��F
N�D��M�����J�v��ES���/��z���EmpnмP��O�Xm/X��jd���MFKgv+Οiڛ�^K�N{\EӉ�*;5N��Ti_�d�
�E���ݜ�Z��>�\��=uP�Կ���f5�,<�K��q(���9�W��8'�*���{N;�>�wb��>�m�ρW�X�4�j��/��i�ݽ�$�V�k�j}�oʞ��n��WM�+��m�.M����V����@��4a�@�fv��6	���0��*��/�|��z��3���YCP�@h���]�cyd?�����;E��rA��3�E��1p���s�����G����� �'�L� ���j ����0�}�x�O��`I�����a�ʿw��B@�U�`�;��ԃL̘�z�����OT�d��%>2Y�m�>ۏ��h*"f\�����x�����5�GH�aS<��{˽��Qd�H[Ţj��OW	vU��������5z�o=&���:`�*�}5z���Z
삥r0W�0�l�D�I�*}�ueT��4��[mI;�	����Uʲ� �FT�(�a�G�iS+��_���! �Z��� )J�)�%?*
ީa��cX�D0��G��r��f��r�*x�&}�>��`ٺ(m��R����}8�`�O�`\��dSLn������pY�]9Q,P9�g�
��~Sy�ls�y����p؋�Ŏn� ���FhC�F$��433��cx|4���YY"��jq�L� 0��a?� _�V�>p���v��݋lv���d2/�����юq���Kb�a��>KܸƆ@-����~RZ����?��&x:I��F��5�^��ES<�|����Үt�:%������
�@�dEY��G���ܜ�]�U�k�p2�k���02��Srk�릢��!|��mYz ���M���Z>Y�jMd���2���L@-O5l|,?�P�G09HB���^�fب���ax�(ٌ�����Ոb��2I�G��ӨƉ��Y�ԁP~���e_Oz2��Ѐ����^�h���ˊ����Q�7jj�h'8C�7�h�������̼l�����٨�7��_�r]O|ǉw�w�*o�s����ߣ���3�4G�Ź��p[��?��g=��%i��Ě0��y����F��
&h=��`����g9��[P�����2N�Rn�	*�ʙ��f��	,F)�a>�XUg4[��PJշ���FY�qvX >#&VS����k��T�<�N�!��ɂ�y.�ubO6�P%:�A)&6���]y��. �}��q<��R�o-E���F���ҟ�>�F���<8|�7 7:9���o�ǰz�,W�ѹ�>k&mQe\J�ѝ��D�ЈcC���6TeL�'g�}[�(\	s�c��"Ȝ�����Uڒ�`��c�y��ʂ{r[t˥̾��&c` �VIL�x���Fh�������2�:m���q�N��R�Ȍ�^B5�1��E�G�~��&}�3��}����Wțe>�V�]��A�/���ˊT}R�J2Z�o��c����[SÏ�b=���=�
�~��}�,�z��f����i�CbnSw���S�������)�e���a��NZ�K�ϤI�E�ĉ�O�)�؊�2��� �xo&��Hހ�:�2���z�غD�lN�m���:,���l�2#R�C�eS�`�����WLJ�d]᫵[U��4i�����QQeY�p9N��"H�-((ݠ`�
J��A��`���%��((��
P�@@�H����
I%�P�(�=�ܺ83��������Y�캧�N�~�ާnյI8��!�A��J����"��~R1I�솜�w�|�b!�����L�D�t���z�L.=YW�3�|����q�O�B͚o{��J����y7ﲛeV��V�1��p�g���]�\[�u��l��jƝ��ؐ�"��>;��R��sb%P{;���6:@�D�>�*|v���Ws����|9�S�fBMz�
g͎������Ǐw����M�FȯKm}���ۙ����b<���[K�e~�l�@��MZ�[�R�B�`]�j�Ǩ�&���aA��5U����"�@o\r���'���|ˋ,_�9�/F@C'�:S��uG�������1�LT���/��б*���NN+�Ӛ��W/"b"L� �aP��Z*��ƀϘ�D��K��1>����m���_�o\��`�ᣩ��"Y��x5� ؄���j7��|��~R���rF�l���`�rwJٛu�)%�W�|fS��e긠M?R���+)\lST��v����xh��.�K��:�s�B'�x�����LVS�cL��|�#	�e�
��WfWz��ښ��di�}�Xaz��˸�AT�X����<\����xY@Y����.����+���f4��Dwd9{�����a����m���<��B�󄴧�gظ��+�/o���MԢs1����R�
�t��v�x��naU(�'#"9�3�=~u"����}#��CQ�C򩣔��"фn��ya_�Q�2�Ⴡ���"�!��:��z����+g롻��vY�J>���9[#$���}rB��}�E�n�F7&�;��+�<u�p�3t��z����%#���j�g�q�R�p�ͳ!�����k�/s��w5���n�io�'z���6���������5fg�К��慬�Z�{҅�4w���/��)�>n�D&�����kG^֏��,����poI�����M�v�?XM�r?��:����4j���jw3�m�m�qeN��zy�4F���U�"0?(���	�s�v<��,l�q 1�)HQ'ݬt}V�t�8�`Ej�_���	�yq�
Œ��= T������4<ߔ�E>+�e��5h:��j���."ty�k���{�qrs���'ݭ<]������0�),����gh�Qn��"
���zw�m��R[���F���*v��8��k������Gr^�D�ls
Wy��y��^Qp�cX�5h�c}�����p���u�����Y��;��9P(�/�)w*�G��1�'���f�H����8�kj��(���i��*�ӏ[z�DLz#4e#��S���@��Ͼ����:]c�Zg�h�0׾D�"�h��z��W��w���R4UN�)�1��i#���Ҁ������CEe��NJ;�0��A�6��E��zW>�\��Z�#mU�&�k��̳�v�fҳ��0^�p�q��lKp��9:���,ȭ8OH#Fπ��U�<㧥��a��S�^yu�F9�2���u�;��F�һۣ� �$6���������͍mor|�{�P�c��3��S��x�b.uc��~-�iq�]�Bd���]�����ՀJT�꼀���pM��pi�'�+/fl��}��l���� ���Qv��-�j�Y�(F�6x�Dz���!�	\��n[�ݓ�%�q=�B��Ḟa��_ ��nμ+^.7[����W�u?��c
�b���c%astPv�7�e��5UgT���'�����,�G���^�ͯϳ?}/�W�B	u�ݸ��M�~2�"�3���]�����	�>�+���sz~�*��2���+����1}:�N�䩛��YgX�̌�`�u�˼@&�{g?�0�����:7��A�Z���bwa2�E�B�ʂj������\��
�a�B�cF������=��=ν��Eh-�ܞ]��M8��t>h��ʼ�њ<��;>�|�X�T�f���h������`��~��צ�L��.�9my��5�'�֠����E�<k\(q�h������w��Jc��_`n��Z�)5['�>���¼�lwƳ�Z��2u����Y�~��1��=�S�ݒQ6�Q�{�0׵=�\'� �[�r<��-�F�5�o��f˟_|%P*���#O�P#����HѴ�ò�����wҰst�W�w�0�E�(�y�W��%�U?����J�Z�]��˅�.wݰ݋������)*�Z,M.|�����m�]��ȓV���*�!%�n
�
���s�P�HF�9>lwxc!�:,�v�}8{{q�FżZ��F��,� ?�L0�ȵ�҇���G�%N��8C���M]�Y�����\qo���8�r�u:���4����X���.�"�6 ���'΢-�����`�T�A M�~�z�U4o)U9���CP�$��3*Sx��YO6Ep����.���7�j�y:��U�+ZT��gTs��|	R�NNЉ�Ivr�є�ީ�4F���eV
�����C�
�%���u��z=^H����C�����Nkj�
����f��aa�g��`�܉�k��:Hq��5�mϰ���	��ڱ�	����!�X� ��:�x��@���ʹn�u4]l	r�xz���o�g��%cx;���.�(�NG�F@��������4�I��tIy�hW��`[>#l��@P#t��&;Y�
j�k�9ۍ��������Zt��`���k����:�D���m:Ʉ�*��̲7�d�6On�P����#T8`�L�j�P�V(�]�#��;�g��aq�SQ���7q;�I�����q\ͭ�Z�~`X>$���6!�m=5�_�2%u����znW����@��e����Z�_K����%�sD��Mn`5NF���I�*v�O���t����)O�z�η�/c�������8����5�������X��-�쇍i���u��M�8%��Ɋ������s<�Π��p�} �,� ��mU�Zâ�  5���6�V�5��("0nElJ���(b꾾�_[��Z���;�ɢR?�C`͡p�SC�92�&:N�D�Z)�,2�AL�b�k��Y0��4a����g�ݐ�5��o-$)�^�GjB�e��Nmw���%�-��IX�.�DL(e�~�����s
>d��&�m9�RpFG�ܼ���|'�iv�Q�B_��C��L�N�_OS�-p�zd������P��`{`�s1�4�9�Qǎ��Ԑ�t�#��c�GF�g'���gG�u��}�<���]^b�=�3��{�����[XwGYz��b/=���I/�t�䡝�"��L}���%i�ߔ}�����Pxw�}��^X����'��E-&C
Ղ5�܅�����dY���.������ݗ��^�oـi!�����Ӗ��\r�;��!.�0����f��|"h�k�����h����\��,s���:��n/vʱ<�k��X\c^6s�m�9��������sH¾��7<,~/�M�� B�ܘ;3�$~�z�M��?l�����;z@ӑ3J�l];Th�>xC#a��g�9�[`k�kZ�<ǹ�N+��}j����k��[���=�,�ry\}p���H���(c���Jx��y<d�wa��I��ɸC��]��Z��o+�ο4�y��d�<�Z{���t<�Nmi'�c	��GU]2�I��Ȥ�����}:�����sA�Ōk��W��Ż�"_|n�����X�6Ӻ�e)�*�
����^2a[�8�P�$E�kh͞}r��Ǚ|qqw��8�ӑ��oP�qz�u�&m�]��-�Ƙ����"��7���R�I�5���y�ft��ΡО���,v?�9Ğ����.�q:��1x�Ξ�/+�1�$@���}����ڧ�B8Xٱ��1�����A���z�`�t��}`�&����84zMa���p�h!�����@9^q��Y2���V���}�@��'4f��>o���@����^��#x2_�AN���RT�e�^4��7a�]i��i�C�{Dx2�|������U��z���	�N��,�N�4��	�:��9Y�umo�ƪ>�w?��	�v�}{j��1Z�!��ׯI�~��P�C��^
z9�|���������)�e.!J�i�)�G�ŉ�X �7* ��a֪ajA������U�<�џZ�߃�a���J�w���/�Ã���5��NKr�Y��>��]���AKz��W'+�Ѻ+;�����c�b��@�~��k�1q�(�|P���1b��'Z�k�:V�;�6������.7� �T.�\4Q"����	�)��J�� ���j��\����]Rh���KĜV���Q=۞�uKiK����D����`��B�=�$Y6�:�)���c>�s$*, ���@����C�[�kc9���3�zP?� ����>IX�Wj?{?3|�n���ʶ���I�D�����e�ƿ�����5
�u�t�;��Y8B�q��Z@;��_n�M�l�B;iHϛ6�g۫� �������S??�����Hf~������\G=���ю�b�)�耲�E_���?��d}i.o0~��C<�̀���s9�/�-����-��K�u��*(>ة�?���k�nv�@�ځ0��u7��p�F[n`������k�_ƃ^k{4.?o-������@����6�1um*�˫�_�M̹Г	S�؎<z��3���r�Z�5�·DLt�DT�꥟c^�i�=m)�"����>0���J,̕�a�+;�ڇ�k%5��M��( S2�����]b��.8����iv�+?�~��NKI���[��}�|-��P~���=������S=y�o�����<F;i!�����n���$dk�u�3w$x�/��Gئ�8��U%����؝f��������h A#2a�O�O�,����=my�����B���M�g�-�?��#-��F�fꎃ�9��3�𖻔=���1+��A8ᑠU7�(���=f��Vg��K2Js�;
>����:��EO����`�fm�vD�t���u��a����x+�iԎ�9)����՛ﻔ�n��0i\7=�$r� ��x8]��v�l�ů���DHw�c�Q*�VW�Xd�1h��s.�(8~�0�ԯM(�tK�Hn&�\Je�_̸�8v3/X��i�_V'ҫ���&	Y����6��ՎNWqe�:-[Kr��lC���#���U�;�:��\g6r���]�,��IX4Z�w�����3�g������Ŀ��{^�.����"�*����!�V�����ڜ��9�%����+�C��xv&�H������yq��\�e��n_�=���]+��6ފn��$k�̭��5L��={�����
�����on�O,�ۗ��O�,֍����w+����sRC��,T1����Gqe�P��ç��x��7�e�W�s�x𾯚$L�D���W������e":P��0_}t���Kk�c�VT�~%����[|+��*-0@O�2z�D�p����>�\���o^�Y�d��_�xsq����^��?[�Yӳ[���)R�������^����+�EG5�UJ�@O��@\]]�^�f�$'g�"��(���D��F���
��7'2c���O�N��{���+���y�����|&	o:��Gχ"6%h���7��]�ǁI���t�ʸ�s0���;�|]�eT]h�h���;0���|i���쎱��r��ݾ6[�������מ���ү��k��7?ؙ�^�zc��Μ���"��:�9V����M������کo�rq��f7븓��եz���~�����dwXk���èSB�)l�h9��a�3Jc�r
7���;�o��w�8������%�z���+{�'���C꩏/���$ǫ�����\+�} �x}:�n��i�?R����������È�=ն�J���ӣ~��Y�+�_��Ƹ�U_;`���.�Jѽ&���n5��U�Gf�,^��L0�5�
��)p]��1A%�+!���k�Y�����7�-�;-���Łm&����LwJC��[#[v����h�R@��߉���R�_��k��u(1�����m�Qe�A`�Wz��1!��U�o�?ޯk�dXx"t��wA�dc9}�A�{�S����@>��*��tDS��b��<e�ɇ�H�]�}[b����8^��op=��4�= �?�9[�b�W��e@�7j�	_,1���K&�9�J�n>�.��<������Q�m
emIl�\7�%�x���f���m�r���͋�*�\��jsk�4������Ot�V5�1,�;��o��x`�-$�/�Ә�F�P��b�7���&�e�%�ŧ>F1�J��,:w�<�O3�� �y�1YQޛ�T������݃�=ѡ���h��f���m�
���M��Z��G�D�ǻ�|W:���{<e`�o��֬��5Y�Mi�/�pe�oc|}}a�N�{��
w9�͢~�+��D|lՄ�hq����G�3�����vsxh=yS�{:�#!��^����vB��E�(����9�R%�����J&��zeG�{�E4+v�Z����;�W�9�>dg�4�˿��9Y��q��l|�N��A�����O*�_��Ϫ�M�Ay���Ŏ��iQ�Į��JW͐2_��D{��{������M�T`f��C��[�S��(���|�Z�r_l,�`�e��53��#W��ROR-���[�Jl<J!���7wl�p�/�n�{5���(�^>����!ioNJD�餢`E���2�՟l�3TD�>Jf��Z�8�#�R��5�4�����0�����'���i�����_���)M�l)������!�j6nes��s=Z��+�3���ٗg�Y�IP�/�y��ce��q���si�������d��RQWN���nU��]�e����¦�����	�����	
[P0���L[�~��	z�����������%wFR�,��Fʍ���O�Άv;1�<A����!=�ۂ�R�I�V�/$�RM��0�Z��^��a��?s�T�K�I�VL�ӑƮ�lf�/B�->�l�/��O�'وN�S�O��Z�N�tS��@��rK�IԣV#fN�L}�$�Q�o��8���yO;]s{�cE�y�X���Rp���rM:���]�n٧f���kb�_�pS�<����j�P~�;e`�3�5�r���V�|/`zG����ϾA=7?�()Y���{��.���[��ݯ���Ӿͫ�I����ܠ�F*���Ƈ&n/�L������Y��Φ�Vz฿�˂����b�b���F9�0��}��5�������Q
c��R�%��E��=��/�t�[�Z��z&L�μ��,�m�ut�>��K�E�9u5=�2C��Ç������Ǆ����
����?d��"�)���o}�_������Zh�������������D>����o"���&��o"���&��o"���&��o"���Md�F����W���[���(s�ƫ��n��s֫l��>�� �rY'�����Đ�z?����IOl�����e���������V����_��&��o�	�&��o�	�&��o�	�*��������o�	�&��c�jW.G|��W'����v�v�&�@�����v
�%�K�(E_&����wyU��k�\m���������(ܾ��8�형�lL�����MtK���/��p���{����ȣ�ˮ��𳔓�/�Ô��WyC���`F*nn�_TT�O��z��EWp�g���
5��̢���G���#��8���Ƿ���7ӡ,��7�-�`�x�~��JB��׷ֽXu���p�C����*'�y˹m��jNӄ�@�Mo%j&7ה�_���[��"A����{�a݆��Ug)�����l��� �ɋ�|imfj�^�ݱ�ɉǺY��}#s��c�˨B����O�XK�Ǻ���U���6�-e��?^�&���h%��o��{QRRr#sS���u3.�k�5q\�Y<��ʲ�X��򔢬ۺ��Q���la~ў0��y�����\�Ù�}��e�w�<�j���gT���	�臢R{�FW�zH�����k~OϾ��w؝�[��X\r����A:䑳�w�)E	K[�>������3�ܧ<��}�@�E"�E��[�X�r���M�w#�Z��N����ػ��3,:� n�8F�f�LK0���$i�F�E9!�c(~�'�W��Kz�hg3�;A�s+k�!!h�ٯۈs�����ϫs���^�(��_7ISeŻi��گ����E՛�	3�.cJ�Xl�?]���DO�@
�9��Η'�eD�1�̾�(�b�������O1�)>-���\|~��(#���8����twKKKg�G�&�~4�\�H��m�Ǧ�{�ĸOHJ.f}Fˤ6��:H�?u��f��f�J��+!�O�����O~�Zز�6��HW,�ʚ2z�6�a��[�����&d���ę\����u R^�7���F���|���+�F����{�5^wY{3(NƁ���w#ΩUUUB�h�)�mX�R�M��_�˾D*4���>����rXU&.d�!(����ۜ%:k��)�*�*G-*C�5mڇ�/N����us̲p�������\]��G��'H]�h\��?e	{��җ\TUUW��AW#��]wumy�/%�t��)؂N-�NY �7w1R<�-�as���D��//�uY�L�Ѽ���T�f��Xu���ER�-w��/OY5M�y��`J��������n�Ͷ�3�e�D�d߂��r�5�S��U[UWW����}�e�y{����u�Dt�����3��Oi;1��%L�������^g�����(`E����`�؛7��m[����i�Y� �#q��Ν;o����A�,��&ƽjR��7�2qm�Z���R'qO�o�������gm� �<�������ϕ+�x0����Z$xq�D#yv95U$ ��[h�O`�WF��Ow�1��p��v��+�:�(�>k�ak�o�3v�8�lp�Ό�rqq�+`��􋰰p�9�.�9�ͷ���=O���n�ދ,z��{���CZ��Ζ����i�q��(+�۳���ʒ������G�1\*�cA'qϽ��=v�#D�T��l`�-{�i�����(����9�G�OJJ2�%�`�Nā�K�L��^���S�|���5�
ПgQU�YN3���}E�Q~ ��(m� 0�9�gb,��n�̒u��]\ḇ��;<&��&ɔm��b$�+J�� �^b�oꞚ��M� �	Fh��W�2'ǣ�#�/�q�)�.fx;��wqD�j�@�m%=� �̯�l�Ǭ]˲^���ƽ�T�VgM��~�yA��=afVzw�����(��e����A��S%y6����O�摈U߹�����D�k������OM��n`���j�U�B'�Kw�l�Nn�I_�x��Һ>H4�*��bۊ�"�2���6�@�:��$�+y7pI��`�k�vQ��.2Y�,�@	Ϸf�c ~9��ɝ�*����#(K"���>�\�돸hPL���C�y6	{P�v��+��ńF��Q�p4R����b�A俬6�/�N�k���A�#�L��VWW��X~0����)tҵ8������L`�L���@��������+�z��'�V/���U�� ﹐BٍT��U	���~A�H"�ވf՘�|i�/S	��0��[i���qUn�ḪaN"D�b�(�Z��"��Y䭱�,��=�� )W��4�.k㘪ś��I� ��x��/��ܹ�d�f\Ov�S��aPf�Å4d0g��Q������k��=�Î�Siii�ǿ�,���?��p�"��	�����}f�fà�,�:�=�o!�}*c��L�g���`���S�#)
�q���x�eӭp�"��}�36i	kU��q�0hmm��I��Z��&�y�0 �����)�����LY�(I6�	h���q�g���VlD�3ov.l� t���R�:�[�)��'Ѧ��"k������d��oġ�$�2b�¶i"�򼔔�s�t���]�Q�%�g]���\aQ|���e��I��&G��)M6���&?!�؋�<2�U����Xg����̩�Y�p�$�_tH�b�d�u��i��O�8*Y&x�T&L���}~077�m~eM��^'6%EGG���Z��kp��v;6�p8�cjΡ��&�R����=�m��:������+B�����!i/�y�J�s��Lp���Y�����d�yv�h'a."�Kn��)�ri� ���C}#�ə��P��xg";^
 W���/���򜄬R۸]v�DZ |g�j�Μ�8��̿tb�d�t�^�dG�Gi��
rHx�S��N���F�(��t��D=h�5n�]�R��S�����eP�g$N����B�2��^ߍq"�7��,yiF4,(����'�TE�n�F8`�ƅi%%�1{�T\�B��e&�z�S�&���ƛ����� m�Xޞ7>��~��.�Z)�62ȔA�2��od���Y29M�!�Ǚ�ϵ�N0|����ݛ%�w#*�ï6|����H��<v?j_!��,΋FN�_�Ci^x9&*���,��=6�*@��d��U�{Oq��ރG=�n����B���ߣ��ֲti�����i\��W���9�'!���n5K�Q@C	9I,�ȅF�}P)?���㛒zt�=t[��c�TY0��fxBL������ǲ,���z⦪��R���T�����ZSSS�g�Tg�X��g%A�蛙�Q'����mc�P�ؽ�Gi҇�1|>��S�$�wR�J(n<{琢��i���x�2V�^�N�,--�`"� ��+��v��+�A�Ӻ��u1�i�.�zK���5З=���� 4��Mi�� %���{OyA�sD<Sx���e�������kݠ�r@I^a�+4h�V����,7ۄ���j*��[����n�6H�g>�u��k�c���7�>��V��:��|/"�J�.2q�4���x��:;n��s��n�����>�|J��y�֌D�La.�"�'��R�	PǸe8�˝��!�
�7���<�H#	H�l�&
Q�vO|��C��6�.J��q�M�F���""͐�[��"���*�n����y�b�Ni�a?��d|3fX[#���&��F�}T\�#Җ�l$��<�j7���ꃲ'�J"����X�Ƣ9���������I�0��͵�Q���~S7V���2B[(W�Rm���m�"Ng�gC��<��]�`Z��v1O8�d�"k�Z��z�)=�PŮ��w� yh0ªk�gS��֎"`n�����y[�W�3W�͇�)M&��
0���~��,*;��Y������VDZ�\4�-�X|i��Y��r#�~++��$��@a.�Ir��|��r#[�!��{/T��N^��ld�h�}tɑ��7���/q(�����d�x\is0��6��)�K2J@7���ㄫs�LN��nwi��A{/������&&姱�I�^g^����%IԴHI��ӳ�ެ�PfB`=�.�27�,I&�������e���J@q�!�Ҟ��^�*6W���V!�@��-�jծ��(T[M���D�!�X�����m����Y��'0�D����g��FCM4��Q����ޗ�>'���ĺ>wo@�b�ߏ8���+b�M�q]��.��X-�٘4r7�f�	S?�b�-��yb)�s���j3�ld�S/<t� uU��)�%L�x�TD3��<�ǒ�Ⳮ��HW��O�L��.��=�ʍ�Q����§i ��LL|W���_#��<0��/��Ҥ�0 ����n��FEDA|�x���JT����u3��4�2&�����r��h�eh�M�z�%�dܹsg2 [�{��ø��J������+E�X�l�
	�(M���G���6hLU@�.\w���T��S�D�n�V��"KS*��q��W^0�8�F���������J:''��)ER�Z�V����fyJj�N�<<:a$�N�-���1K�3�o�`i�z�s�����m�����*}�6�]id\5>M |:�g�'WR�j���X��aZ�uO�Կ%�(����У��4�NBz�3��\; w�^����9���ݩ3O�\�8b���������%����;�t�@�e��2?>>�?Q'-
����U�8��$��˗�	�'1vbܫ$��$<�S����6�Gp_6��O)�+�gK��gH����0���;���c���&���R��OP:n�}�۵��'����kl�,��
O*v{*�F�\�6n`W����_� �w�2BQC^�������	l�T�x�΅��Ԓ��p0��fC�Ջ��3"�$`�̑Dq|���FǕ�����PR�T#����BZ�to�Q~Ď�dބ�4a�?:�2s ����6�B*Lbx~,N�ӕH��By��D�!�>�vۍ��ٗ�-7I#Ch��3JS��j�6�N�ҷng_����ݒ4�'&I;���ke��㠡&�� Ȃ�巐���@��/��07���F&`T��xc��}��d.,�qw� �Dժ��<����e�!�ۅq�Jh�ܐJ�򇩓�x}�+5e��7�6m�m(���&S�O�c9���8'���A���z/ GO���`!���\x��? ����sƨ�����D�?��W���8����d�Y�
����8��Q m�j��`ⵇh�nnn�K�������^�slhӗj��,�XIM�Xn�V�T��p��:����q���ڬ"����\vƟ�;J�҂���q�6:�y�������>���"���d�/�$J���W�V츭Z�B����Z��\�BT�e`�Mc����(-c>��ێ���I��7��o�\�^�+�ku�!�k{`rr�]|BBB
g�'�3��d�)3k�C���o`�8��J�y�����P�ո/c��_��@@E�L�F�U�/(+��5j�8�|AgK-� Y�4	��á����tn�����:y&�W��IQ��C���n�$��LC�6�+�}&���c���6H�cO@�yaÌ��\8���S�ƦqW���^K��'CCC���rK�_�Y����+=s�҄��<�Vttu'�;v`r3q��ϟ?71�����+��<��Kr
�j�%�s��C��Aǐ����y�$s��!������K	D�j�휩�-��(TX�:�U[�e�@���U�Fh��z�VE��{�@ ؏f�Ct�%[����?֑��A�>��+�(:2�����\��=IM�-�y)�Ҵ��s�$&6Vv7X� J~NR��o�"�2B�/�5�2%%��8�@��q��K���B~�\����%�6�?����b�%��i�0\����h�,������(-q`��o/�Ft?�Q�� yj�B��C[[{�0mN�u�V�f���&�V�[qs�?�z'�I>�m��ӟ0�\�Ч��KN��d�n�ֻ���㜜���$���w;�{�YFT����7���C7h����Nt	y0`�����U'�&o�cw�^Pwʓ)���k�͑�p�8�醟y��P����Cm���@C+]�z��Q���h��k0muK3� ��%���e|+�2����=�Η%%�M`��>a�Ά�m�-���3��@V�`��b���y� �%��2cz>jB��G�`��Aט_GG���R�ص�"���](�W���U�_60X)�4�A��/��f����%��Φ�[���\#%��}���4C��C�|�t;�zz�Z6��쮕f�$���.~<?������I\#�uy8d����h����e`���g^� �=�ow���z�о�y��U}}}:k�d�,� �[���鑰��E>�tL´�r�"�>��.�x���3Z$Q�ç��z�$��iw#.���D;QZ�Q���{腧�(��N���M�6�?ͻk(��ێ�O�C��~�� R��~
&`�*���DE˽mm'������(l|�w�V�$�&�bb����_�;<Y	0[m-)Bk�R0�����gձ���	�1ץ��+�� ����ˎ��z�GH�Gz ����.��\ns_��u��cD���k�-ΟQ=����e1��w�_��4���+���jN�&����n��ݿҷ���Ͽ�#�I�q��gǘ[�6J]��:���o����w��=־�䛜t��@�XI���ť�g�tn�5(\fb�%/��B�0O��0Vx�?CB\�#gv�e�0�(�\|h��VIՌ����(���<�}�����b����p�k��/�����qq~�87VXX��:���}���b���;��J� ��=>�������A��$U�ʇG���g9�ui@��wk�t�l�8D�w�����LΕ��ù�
�+�q�@��5��L Ns�@�$<�ʜ�9��{3U!"����%�e�_'п��1;J���i��Ũ��ַ��h�G���R^�J^�`n�(��.�`$���:=D(��S:�=Ϧ��l�*	B��M~�832*j�"ʚN���ƙ���YaU���2W_r�={��H���v�����I	�`Ȇ'�y�7L�͇����q��>���[�'�tpN�4&2��UN|�����D�Fg��f����5RM!R�A��٦g�f#K�Lvq�������K�ž�v�ymT�6c=�Sj��
�P�jhl,��`�FA��8��\��I���ir&�G�f\ll�����Rt�����4]��T1 �64�bk���qa2�9k�٣��4mR&:巉N�|En�����v����DvQQ�4�z��?����N�R�nL\7�.�u7$<\��ral�)}a����C�t�l��G(M�Q���b㔦�ؤ�V�I�b?�*v0i,P�8T�ґ+i�n?_[[G�#�~C	�P���V&P�vD�E�r"s��Wn��>*�r���K�?�Tys�뎹,�l��W}�Q����Ck��b����r��\_��vS�/�!͕�:=2��~�.���b@ ���N��7S}��=�MH(?¯�����P��EP\���n�5>m���Q���R�"(���x�-�f	�a��7<��c��t+|�$EVΪ�Rg�_�N-w�%hABټi��ߟ�(� m'X�Ej422*����C���eY"x�L�U�d"�8Y\�� jN4J��s(��:i�K�VM�I�Z�nr9/w��Zrs񔕼R �]l��R� �-W1P�ow|`ίk*�	�߅Y/��Tt%��?X�}x��xr+�E���H36:&�H$~�AP��e���yү$����Aۼr��=�h������@j���A��YZZb����� �j^�'�/A_R,�r�1,�.��/�!���� ObX\^/�(����@SX�.��	��ﱵA��\�y����6OT��p$�]��f,F@���lr���7#-۾��)��Հ/�0�ڃ(M� Y&G!�g������u�̍��Eg�9�Х������/^5l�;2q�|�t��,:�ejl���Q[2���9	��" x��;�'$%���L�m`Zy��]�u�K�C<...���U�|�#諹����C��?�X����j����62�}X(W�D��}Q��} ����CU�2�
�Eb�Џ�!y8Ya�@���t0VbC��X[��{J��
�Z�X?��y�6�J_�B���]	u's�t,kG��^J	r����2��2J
-c$�zJW((ӄbYId/�qU�j�w��ƺ
gE����I����ׇG���h�U�Do�FRDDĤ�����s��"E��_'+W� ,�� ���zʁ�`_��҅٪X#m��3[�0XWW��Jj�~WkHjjj�J%��e�9���޼�\��7:�6����V��K3�Wָ�J�\~f$␶���w�f(E$õ< ���D�o4�D�7���Ci�����ح�(ÂG}^|ޫ� ��&ps���U���g=]XX�3�7:�<���y3�G�*��U��+D�]���B���
@�%Q�W���ǰ�E�H�.[�/4�ɓ��Q��_���v��^����q?*�se�{�9Hr�nNN�������h��(���2�f5bi)����ӡ�:�-���=�:�'t��b�ER����&+)��4�w�<-�����J������4��6(	~�K�z'�0�xV�|��0��ߩy/�W��)����lx�-7�)��W�CNA����[�J^�M��z�7:A���{�� e$���"�	e"�U*�e�`/��Ao@y���R"��p�}�s���U���Z1�z�~����lC�ߘH���<q͞42�a%
���\���K�*ʃ��/��!Q�Y�6��H�����r�btt4��P#��b��Vu�	��>S����B���6b�|��E�n��V����ٶ5"�M��(ߓ���[+������J���� ѐ�ds�=�En���O�R����=N�M�j	���a��L�"��` ���3�l^���q[��В��~�Z* �߉�8�H��_+m"�R�6�@������ݒ("���H�&�-����@8��{=����{��0O�,�ۂ�KFAI�O.��#�}�y���t0�|�	��cz�}��z��Aj������bo�f	�c�}j�����ݹs�SO�gch �c{�E�to�DG$�*��K54j˯��@3�Y�L_�$ю�^�)��NC������%%�<����A<rj�-��p�P|	b�\�ٶ/K#8@��Y,��de��4*Uj�T�#����^�����sYд����͹�NL���3uĩ��<(ȏ��(�U�𮯡ۇ��%���f�T"��T��?[ZZ�ӟ?�B!���0��Y���@e~�����8Y�Zֳ�,355�s�
2�T�
�-�pY:Z�ϐ~��@�f@wg�v~^� h�<�Gg��K�e��T�8��y���S�L�E|!��v�~�2i-7�A�p��\�KLg�޽w�x-�ȟAЬ���i�B��"�J6��*�S����ZE���ǥVQQQ|�h%�R/��l��+55;X�K< ㋷�~���:&0�<��/�n��d�_�)(�-�J%)�1\H�V�l���MO�R`�����h!Y�������|#� �������^��JK�E�%���n�Y��f�A.Nd��!j��m�u?��g��� mHP�H���f�eA���i�[g���Ql��S��G�do9��\@J����뻻�>:1R`��7����R`��^Na$�F�/��X�����N#ᴸ'�LBw+�C*I�6f*��R>:����G��S�H ����������<k�^�nb�:����S�ՊW���Y��ô�u�ʴ��QJS ��KCf���$T	`h4�[?L�:w��T&������#�����
���fdNy���)W^�\�:x�H�'��Ǣ��B/��{�&Q�`���&�gym�5�~�'�z}����5�����p��O�����lT�^��ߓ���̿s��˷Z:�L��4"V�W�Ł~ о����UG�1؄T��S{����N��J�Ԫ�]��'�@酻*�؊q����?�'hO�,F)W��Zn���9=��4K����)��#YvL�0����V��%�C��y�g���ǝ��� �XE��suz!�]Q8�~=V"lh�mo�a>�$�� ��m[�hQޝ-����;��)�cǎ�I�v����p+!(<���P�>��i��n���s�N�V��pJ���.�$�@v)�"U�����!�1��?rf��5L4y��@Q�p�"n~l*\p�[iEx,z ?��<X"�\�;v�rp�f/�y�T��O{�����u��)+=|`�;u��H�9�E����ǈ��̋�6���1Gz������z���as��B1d.SWGgBj+��$+�?����T�������|;�R��[���˃��X����#}���u���W}��6O���5���3�C#r�����(E�Y�5��vpY�&i���OS�+R��w,������6��g�\��4�R��)��Ν;_����X�C�u���ʒǎ�N���S��a����@u0����P#�6�oB,�Qi�o�4 xu-�f�T�Q�hOQ��L��~#�ߞ�i����3,\����]-��&S}\Q�Ͻ܅Z���haG4�~HS����Y����f�eܜu�Im%i1�©���9�RiF #��ã�Ux��&���2�@�^�
�y{@T	�7C����>�#ӆ	���<l�z ����ܢ�9��N�[�'���=��R�8̿�Bf������(��
|�?9[�7J���j�T�3?;F&tnv�	h,�/�[��%��� q��;�;�<\#���QH�'N���36.3���Q����v�NUL+�t�:h�f�\���.S~�"��A�]�[��g6�FG`�#�'m@���}󺛑F^˺�����ss�Zr���U�c��@;]?YV���p�(/�X��� ��'�ɐɃ�*��9��@y�9���iu�Z'm���5< �٠0��a��@&jb���D��X��$��yo������1�s\E�2!
��~v>H1_��Mَ������rN'c�Ϲ���v��b� ����D6<hx�9�ďM�k�T������TL^�����|����ن�C��/{o���B3��
)|:�'������R(M�T�7,!�@�Dy�ܤ6�%�m:��\���,]��Q�;��z�|$�4Z�Sy��?��v刃�ٖa��i)NI�f�Q@��7���
Ӓ��x��)����~Z�j�:0�*��6Ee*�AAQqG�
deY�DA��j�4aɰ��(� K�,���w�r�������3�w��C_ov��1j����F�7���?4�J!E�
�^ǣCW����!�Ą�ҹR�/�k,8��o=G�[J��	��3����)�3}���}fUku��M_�p|\��=�%u,�c]Gkkk9�����AR�/ى��Q�MaRRXVRVfq_��n��Dg���anV:p#��w���e�M��Ōҋ\U�#z�\zh��Ǒ��=����g=���5P�l������	�g({�:�s�T_PA�Z��Bk����dp�����|wq!��Ǧ�#��5�?N�IS�8��0�Xy��{���\��s�[�g5�^⠅��6nV�jv�mX�(�x���\���#�������ǙuO@�WY���t�����e�n�f�� Eދ;>��K�y�C��� ��*'��s���P��E}�VnZ�5ZI��fY�s޻wo�@������}�?`:9ސ��t�޽�cy��I���?�s)��ܺt��/e����x��/\͝hD��9uy�����l��Ӟ�n{[���&SZ�s�����ㅀ��S�}6Z�!L��t`��t�vIFg4� , ��;��!@�:���r=2��xK��)3e#��i��ɂ�.�u|m1;;��4d䩅��+F����^3<6�������傕�5io��G���b�r(`�j	��Q��L�5Y���w���x��}�&¸t�̕���줾��] aT`p.=gc���vP�i�z�ܹ�{��>Ҳ0���Mj�ճ8��;ǜ={<�ѿ�����^h5'�ɚT�GsȀ�I��]�6U�Wj�����R�{wd/��<�@�G��g+�b6��*���o޼�B���V����" �X�y?źf�Kt+�f���>���т���w�)���K��#�u��8ٵ�<3Ea�.c4��[1d�|����U�cGM<�L��������n[mq���K�c�x�N��/h�=�I�P_�F*A����^�;d��f�MH��Iofһ��Z5?��3��_vLA�<�>{}u���%�θ�k�Wo����a�f%$h3�,�-Gx�P^���+D��#�^�w�Y��^*&"����TR�Ϳ$�n�u�3���P����F��K=�0��l���2:ԛ�M1�Ը��P���y ���0���֞�~<ߟǷ \�x�9C#������v�in%�?��ry<[�Zv�H�:2��?"���>Wa���qH������_��.![��٘0mu9}��]9��l^� � T�;a`�t+�t�l�B�s$��ߨq%�粓�<VR�vU���q6ױj�������[{��1שJ	�"H���1f�2�-�dXE�{C���	��򢷇��S�qZ0�ʺn��		
���:*� J�i]:`&�l���e�{W�1����?�]-\����Nj�Ff�C �*�`y0N�D�����nb]}L���hŀs�@*��:���߄�5}n%�v^��f�#j���B��}ł��ʲ]��1u����u/�&" �Kr"��Oѱ����<�=�fy��F��\�)����e��z���]Kv,�#��d_��`��
��,`�&J��8�߭�g�?��ӈ����B��^S}޿�j�,��$M�ka�S{���m�u�=�@�M�Z��4����)N[�\���F�%��}� �:��l���@�t�: ʤ��a�H��0��_��,܋aC6,X�[-�+��p�O�l�6�.<@�#me�IHxϭ�O���h��9@���ѐ��2Cn�Y����b�!gT;�P}��dY꽒�����.�~%�%i� u��TQ�~l[6�Y� ���GaŒ�{�����
�Gv�Q��mY�<���T�{)e�A����n���MK���nX\	��w���f�MZ��޽�4j���utܵ��/;��MG��Ka���>W�o��B?�ҭV_�.9����?M-޼��}�Ϝ��W[_�:k��)k���s+����By�[��۶�¬�?���l��fz� o���7|�����|Y��*nȻwʮ�׫�v��<~�5W�ox�CB�Z\i[[��D����|�f(��j�P�6��*Ca�&�*ԫ����ȍLG�l��4���[�y��־�	���/Ճ�c��|>�~d�s���J��X^dN�b��s���0!��P�HYc޼y��!j�� ����Q_f��QZ��]qs���ن�����f���Xu�ج�*⪪����^���d^s�ݳ�ɥ����2��6yp�nvke����'�����U�r�8�gb+�a���D]m����13739��:�8K��ϒ^7��.��9 ���5���#;�!���t���?����,omjXɴ����I���@-2�X�qʝ�� ś��k}����
�Z�^�\r��ms�^^jjW
�U'����Q�Za���ɸYI���U��s�����hů�~H�;H�������ޡ�pt4&�}C����+AS72�}.��B�ǭ�R
����c �^;PYӌ7U������DJ��F��G�k2�����ϐr�[f��t�1$�y&��>��S@�be�����ݟ�*S��:�fGj{5��Ǐc�mթ���&O�AH~(//_���#{�)璲�'��IN�[˘a����S��0���!��G�����|������] zl(+�ml���@sP�?�ĭV�?��ƄS���=��Fx���g���D_T����)L��r7��X��<i�-X��X���X� ��j���:��Xpa]�C��t#�����i�'���~yx�#\:�|}G��6��5�k�ɓ'W(#N'�n#B\�M����2m�z�ii�1E�el��~@"�0��������ξc��vWG(��Y���ř��7�%sY�Q��UX�?g�(��6�Uc���{ۈ��&�v,�u�%�����b"��&_/{482������3b��f&
F��\����w�%����P�����6>��%+�z~�,�$١Ƙ3g�z�	SXk�v��z�wO���8�"�Zq�~3�ʹ 2J��'��r�X�%w;-��P�6e+5����>���Tzk~�޽�0Ʋ�@iA���K�g҇����bw��\p��?�j��Q�d���+L�s|lǳ�m��}��R-s�[񈾩Dx���c}(���Gg='M���'�̭?e��(}��<�=ɷ�τ�z�|���=�Q�^gѓ��ȢR<�|r����~�X�Xga���6�N���U�X����V̍�b'cQ��]�w��1l���A>
W��+���1Vw)#�"&(��j���Ȍ<V1ŝ}��s7��S�l��u�SQQi��!�!W�^rH'��r�lʄ����l#TfLv�G[�Z����B�	ǽ��s~�����4�Y��d������&�j�n6	!�?�q�ܹ!1��8X�^�>q��! �2�kb��D<��0n`��V�6'�����O"4�w�q5�p��o�7V-���d��q^>��_��W����ɹ�/8���e)[g�k��q��]�x�bU%e����nL<چh����Y�s��m��|��3���s��5���`e_�� R]�(ɰ���5�����x�s��u�L|9j�m��k�ǭ��5"��^�Z��ו�V��E�h�/��>E5w��}/�5��. �B�j6�Eg��\���/WwՈ�))��Ʌ���?�Q>�E)+[��
cR��?>�zZ��n˱ts��0��F�r�X,�RS�YN�Jl-��G�=k���1���K�c?'W�:��yO��%�c���V|ށZ �1f�/N��x��8���L�q��3_(>y�孅&��3�u��SBe7�h�{�%y�������"tkx2N{d~(��sR��=G��ID�v�4�r�����lǗ昃\���Bz~L�:˖_���T���*'�[���$�C�����eDEJc郗�b�}��$���#�W<���k�XB� ����`�K����^�.����Q:���M�[�&�T�,�����~���U[o������Yqqq:'y����ku�	�2���=#�)z��l"!�"*�O`\oqnΪ�:�۸��Y�����@O�����+11��1�	4���B+ԧ�S��֬×Ń�f,��`#wvivY@(�F�c��z�/�xs:h&Ke�ps���$���e����>F���B)0Dq��atC����F�"K]YK\)I�j�Id�MW�l���7�*������_X�nxx�!"/��=��K���f��[��6l
�6�q���Jɷ8ڤ����o�Va�G�r+�r}��=�M���,�i����
��Ul����A ��l��Pl�g+4���9_ӁX�B�$v}�ZG9��Y5�hk���2��N�L�n~�=`�F����\J����e4�S3��9����D����8��4
R��֥\�������q�T@ů(&[�̖Bo��^�P�ۀA�O69�V�v6�]c�*1�"p��ڐQk�����%��hA<�}���E����L�h��@��0,꾥����+&��� ���u&L��$K�b�B'�%'"X
�oː��`<�!�T���W��u�A+�	B��<b]�d��VF�Az�e���-Jr���jʼ爪s�	��o�?oE���9�)?A��_�4v� �w�jߤH���c�X�q�\"�?�
:=$X�u�]���1���1�%�r��.{�H�-��w:�P�b�-�ލ7���/.���ת�M9�U��=gR�
1�cm�sZ��"?%T����D����rO,�(��,�z�h7����"	�MA%�����M�=����oH���t'MpZ�z��w=NH&��N�ژq���O�ѳ��ϯ��ɩ�O?��ƛ2x���^&#7QI�B_�4Xss��A/�@c�'M���c��5(��E4�*_����/����jb�:�7o���*6��5uZ�9߂�cʚ�X�y2�ܥd�GYǄ��i"�5c,�9zכ�_!_���[�Զ���?A��d����F��x�gr=��?�Q4)��.�V	����ty�)Z=e6��*=����V`�1��� ��)P�@�z�-��.ct=.��2�ɓ"Ui�7�ڤch�[
NOҘ���%���d�t����u��h�� -���b�#�wd��U��M�x��XA�ܓ�]��75�ɜ5셾�*��>��Fx��|B�ƂӪU�@n�k����h�Ն嘠:$AY,h����W�M(��C3���-	�ύ��'%'[̒������$>��*���x��@��퇥�qm�:�p�2�hy%R�[@�:��F�[c�J*P�ʔ�e��3������(!.dܘMO��f��h\�`9��4���	ǧ�������|�;D4D�.�st�����M���I�r�ZO��H��m�33�m��H1�ܸ��^�x0�[����J ��X5T����_�K�gүnuQku_�5����>W/�4b[���F�3�̝|��vE@]�qՍ7�7�=0)���e����c�*�t��<���^:jz����y�k��bo��W>����/w(79�S�C`ͤ�������56����������=!K�x���Z�w�o�L�~����P��hR<�i��Q��F|+,�믿b6�N rU��f�4E�c@D���P�R�]��L�	u�q��j�ف���ٳ�]8�d%�b��4;�wS���Q)ӡͯohwW��c�^��f�=��感sQ!�I���������������R6�������_Ϡ}�_�M_�1�Xԏ�o�ba{ �	z��(� �$)A��7[vlCK�7�����G�TVV~ĺn|�h?c��Z�sv�ЗN$�)*Z@+�.���*ӏ)8���;�<�y� 	o���@�6�O��>�%%3����&���ك�c����$�������U��
�FXJ#��r$����|�
_u�Q�Q1;9'+�ݝF��o�P���(�����2�|�U�'05��遁�J��P��照\\>��0�˳���U3���d(Gs�y�P�g� %Hq���$��Zn�\��!�!���v��Vj�`x�͟�4�n���d73V������i��j7`�h���.iZR� ��
���H�mA)B��u�g�r�= ���C5�i���,E˗->��k����Ѱ��'�bhG1�*٪��dܙ=�9�7m��E�?Kz�����N����cyFaaa���$���z%���  R�J�\���`1.A,E����飉�5d^��@�wQA�[����8=��ö�9�u9}Kq����p���f4� ϗ�� �|����y�UW�#Vg�&����;ȗH��5M���Eˇ�7�&?ߥ���%�8��PJO]�~���W�\H�-�2u���78��N4���fՊ����ki|��8GU׻�Q�0&R̎��X�0G1��C���.� ��JVp������9���pw|��9$y�7�-����|�X��`E=�8�"��>9��j0�,�Ӛ%��@>���A�Y��-%++�&��I��fn�,�A�A��rٓ�%�J2	��a5uS���Ji��h�Ϳ�d�� "��`]�xJ��2-7�ŉjkk�}�ҋޅu��N�ڙ��P����qf �#�����=������
]�N>ٶ䪡 ��W�&l�ީ��f�ٔ\�t���
;Ŗ��$��ݑ��}�gZ �i�D跋�s�U��s�Фxu��O��������\Z����{nC?]�ZO���Qs�i9�Gc7�'���$�L�#�����e�޲�S�g�}ǣr�@�rr�
zY�%�Z3��8dk�C��[��E>,WU��wb�~�N&�#^��o�u횗>kx+Z����޾�> b�kB)uL}�<��Ј���I�N�/�		�6��^x�;�#u��CG�{���3�-!�:�P�Q��|���P�������[(�*"�c$^G�1��q� ����Pw������?RRtv������Pr6F�\ �D�� �w�c��%=l�u��U�q|�YӰ*�^=J�>�%�h��}�@��)Q<x��C�����_s�2 ���s�|=MxLn4�s=}p���ӈ:�=rlI3�ʌn���Ŏ��M����I:Zo�|X����0+�ˉuOr�S�M�����z���t�!��.��.�����b?"�-�I��i��q��	�qTS�]���F,cw:�T�2��Q/tV�vq@#���V�
�5B���j-�7�ɚ���}C~3�����?O� |)���7Ѐ��{����y� �����/3`�{)~�A�儘2�y,O���r�${E��[W0h�U߁����x}v����g�(�n��&��\�`���jw��i@x݄�"�Z��cT��J��j.'�k�
�������Ƚ� '�}���<R��{�U?�u�@T��K�����(L�\�]�+�٬ex%��؈�Ox�4���s���,/���KӫG$��7�m<��Xڰ���8�P�����D�KG �۪S��D�ϡDI��%�y)ѹ����⌀���zW!��٭���z�XT	��!s�y�M��0�����\`���^U�A��5�-#~���0� ����y���K�q�oA��?��j� `���Q�J�@�A��1<7d
*Zt�2F�����c�d���ʠ�n
lNms��6'�UԚ:uj��;��d�{���G����_�q�e\�a0���-?d!��cµ�z���C�|=ߨ�k�o
bL�^��T��kwo8���rQ���_��0)��-���b[�BM.E=T�g��W2��!N�]�y�&�PF�'���	�yO�YQ����\�L��|����nj��f١�K�x��u�Q����ܔ P�����΄�� b��l��x8ڦ(L�tj��^j�����pQ�����=��#@���Y˅�n�d�vv�?0�G�J�y/=)1�b�2c~�m��k>�;bbߝi&E��?���Bk�(X������#���]�Q��u���߬G����sKp�{�ă�8D\��S�)����>V��f}�k+��-s��#PC?���c�#1�X�T^� Рq�r�<Iϗw�5���`��=�s���_�D�pM@�}�;�;����B�U��{�%��% \ރMixنl��"����֯c��B�7_���
-(�������C�$������X%b�!Sa���E��>�a?�I�"��th�jh�Z)>g����紧,Ƕ��(0��|I�ҙ�z��uV�7~s����nfZ]����3Sܸ�����=Z����1������;�K�҇����k#}răg�������]�0v�%�zI����X��&��X�&>��h��p=�t�0I|r��6yT�j� 9�R`�Đ�g�A�=��[O���gCX�9�ܖ��<0����r�z�:h�����X�x��%!���I�KC�Н��O����,�q{|�~�&;�i��g�+��\o���2|��j[�Pd*��$�$��80���?�
�ί�H�'���W2�Q��Z���>(��s&�p8�6C�&d�A[�45��CeZF�4�^���\���e��a!H!�4l�z"=-�A��$#��?�j�,S�`�|ve³��B�i-�����A,��3�M��o�mV� ���J��V�Q"�q��zL��������/I�������
]E:��[F/���!2a�ؑ�G_	����CPR��1��'�2 �7��H)D	�&����G_$��`�;�wX��? �6fP��L8���*����������G�����Hv�Ü$� �ig�62��{@��,��@�}����<�������[u-�R��Lg�����6�|��w٭-]�$���Jzc�,Z�7�'Bܛ0�Roo�� �\�`���8F/�6��MUn#GR=1�K |�8jc�����P8:�� 5��;�+�g��yCW�~.��18��XҚ�p����苮@�8�F(q�Y��BSz
��qC_����766����]V�����a&�Ka����"W@�qiii���}�OU�%W���聀���"# *hqޣ���kt'����a=�<�Q��u���~{|>w�Y�L�!��E=&œ�Nx��x����:^b�(�͕
�\���AZF��b�y1�i���cJR�qKvR��j���Zu�eh7R%h?����9/F�7V�+�8L��H+X,���J�u;��x�DQ�h�y̬��˝�ܴ@��;6L,� )_�״U	��4E�y}����gF�@����6	"��h˶R6W
��Φ=����eR���(kV}Ύ���zտ��hjz.c�^�M:��5�G��Ϡ��@͂"��_����6(NЧ�|[�~>=����,���J�~?�z�N~�	���)�͊���>º��ݤß�r�4J+��U�LE���Ķn��i�x@a��E�U��ڿ�rl����a̐e�F��iP*s���Z��ߨ-_�Y�č?]n�ә�I9��s- 7��ʊ+�_���K��9S�[(�?�I����5p��S�Xd�Y󯉵�_Y�ڀo�5�&qBޥ[Z�]�vt�a�ŭ��~Ox����b��åf0/�ا���p6��[�a|�� �Ԏ�XS�	�f-+!���dO���R$�m�[��:��XުG���*�J,�W=�!���A{g���]�-�K:6�F���Q�?���������c8�����Ol|�3�����!��3Q[��bd��
�Kp���Ƭ��Y��PK   ���X��g  n  /   images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.png�xUP�u��{�;�)�AZ����C�I)�-����8��P��+�{���tw��Μ93�pfv�,B��*�  ԠJ��&��q��un���j�	 0�����z�Hj/�w^z��^�V6 ___>GOk+7>W��S) ��AMI^�/�$���Ġu����������1�6�b���w ����(:��9�A�B`hz/�抉���T�K����%U�0�2!54����+|������#�lI�)���ŶE��V�c����m+�h�@.�����9UF�*o�@��Qt&��t�t�DA:2�L��K�H�e0�j8"0��h�����A�a��/�b�V�D�o��휞�H���l	}� }L�~���>��t����|f?�Y�����0)�){��`��o5����1�䩩��-��&�{�6�P��54v�J*c�?Ν/�yޣ���;_�����WF��� �z����ܻ���1)�?�n��9[��j��U�Ҫ|[;9�K:�D"�m�R����7 쟟[�ެ�68��<Sic�"�lM��ljn6b:m�&L��}�pj�������\����ֶJ�U5�tޢL���n�l�)�ox;nx�TY �J��y�I�@��y?E�ʯ���zZ�Ҍ�w�;��T)�?'Q�63�������W��:�@��e���4�R�I`��V��ʿ׋[��^��FS��'kc��������k����$C��7HY�T���H�"n���v+k)6���2�& �gg���;�>=�y������SAJP��f,����ׯZ�:஀[�?�q���Ǚ�UGtY
~s��^�F)O�\��Ý.�`{��3��b�$�[��H�:/7(���D��Y4�zV����;�r�w�Jtw��t��iYuI��>~ɺ��%�^4%����o}�͊��!b���k����PP�N�˺���y^�i���	?	�<��횇
���<疗9ϺN�s���Y�S�nF��r4J[���松>���]!faU����3�:ːG�q_�
���?�君���g��fٮ��v*�	���P�������)��Wic1�&��
�*�QB�#}�,���Jt��Ut6�c�Y�RY����m7�dgF����w�9f`z~���������4�)�n2~��m������遡`W���g'�x���!���+�y��Dx���/ǚ솎q��0�ط��S�<�+�/@� J��,jnn6�FB�YW�1�z���0i��,[����zUiQ;�D���ϽL���HN[��|o�����\m���UU����@�Q�������g�3Y@�/���Xޏ�w;�s�n�%߷�WtMfI�0�c�IUr�{��K�����a�u:S�a�n|�IY��ARĈՈ�:� ����;4�JMP�64���g �6\]a~��u��E��5M�e)����N;�Y���@̬�{V��ɫd}<,�� rp��!wL]ה��V��`�|��L&�E��LJSKy� ��V�;/�w#����(�.��o�L*��P�,���L��f���n*��/f����k�M��C�I��V�{��f�9��e��x�Wڜ{A���S�z�}������:L��3�DR���5s���l��x9�o!�b��9�!��9�����ӖJ#v�2w48SݷwӤ�Y��VL�kR��NX�I��w�L��/�����}��ͧ���^��hx��x��|Ԗ�+�鳵�	��H|:Cu��*Z��j?|8c�{�|N�1)���.LCCSu����L���(���(]�:��@-�/!�7�?�X��M�-�p�.Jjߺ$�s/ls͂��Eg��L�8�:�?���{t	)�|��V�~ܟ�����n��Lu	�gAOB�����Դ��>
�g���xԂ屙�WȖ ��#�!��{�8ğ]�7�F�G}^���8�xڎV+/��f�}�X��}�,�<cj{h,j���~f��gi��Z�陟�`�c@�3��8���`̂܇�7�7+R)wQ6����"z���:�*��F��7�|l���nI�o;u	%�_�ۛ�?>܃�Ѩ&~�	 ��:#K��6
n�F���4epftg��(���Қe��M�o�#�a��%�:$�O(���SH\'dn��DN�O�)�Y��"<����?c�Ǫ���	Y��;���ª;�lH(�)x[t"�"G��<��㬖�r®�k0�&�`��C.�"0��<e���a��@�^�c��",N<�s�9q x���f�\WOL�F����j�&l�f� �����0����=�����	�@L�6Y�Ed��Cy]���N��5?'?_���Y�q|N!u�ʜ�s��u�N`}���$~��g��^�z�qr	J^b�e�T���ouVT6 R �zynZ�e���ۅ(�0���ȗ�<Y�/�hm�K6`ϓ'�L4a4��{�щO����������"�M��8�;>������m+2/�O������2xS_:x���S���P��A$�޳�l�ϞY�(���5��l���M�'ק*������w�}�����Zq(㪯��ϣ�,�݄1��-����E�w�>�k�O��$ܗC�@x�j�]��O��'N�TY���"\���Q��K�iJ�y��1��欎|��q��b�ӽ�#W��T�Q��ݪ�6�E�#g}v�\|)&�Π��!��S�y���k��i�$��f�*����˫"T]P2 Ȧ��$-t8�j�QG �7��XV��#�{��L�v�&g|�|�;I�Q+>T�f�b�+��s.�	�]t�ۃ�cm]N�û8��z���׈0=XX���8l����=�]��x9��^$9�m��r��/���Ɗ(Nwn��X���Ea��z/�ejǫy&�G�A�1��u^�U���e�Rv��	A���L$��t���k󴊧b`�x�`�`m�c�[m|�q����%�`���tl&i��{CwC�W���v��3zB��/�0
�}���j�FχY�e��QeUNh/�e�违:����y��',�[`�Є���l�#�w�-ܳ�ע�yRx�DE�����.B��l<զ�	�b(Ι�O���5i�K��Վ���R�'C�2��Ut��v���R-�U���H��Sh��W�\h�a3Kf"!N�PyMlOB��	��ɦ��T~��p����&��.��`�|S�����YP�H9B��7���'67���!�2RT��l�K>P�����F۞)/���� y�I���I� ݺ�
혷7������v���4��YH��V~8�(�y�E�l#� ߄ϲ�̲�'7@�eV�M �:P�����D���U9&��*(h���p��`�V������Z��ڎ@����Wu���T�xhT� � �ɣ����w|��n�X����7��`���PI�l�� ���}�wd��.�Dj�z�P�1�sB���E�!w���Q�(�����z�Y���H��-S+����D�Gb1N;h	���4A���	��73o��Z/	[)*�PV�"6ӱ1S�$RϠV�+��_��A�>��2;DU�l��
r'F����m��;d�7V�+�YW�H����4��5K�/���z:©��/ؐ�O��n�w���f�eD��<}�?�Ҽ��_)��dz����"��Y(v�+cZ%,�`�UH��(4���ٯ�P�e�+�靑A*&�4Xf�%�#��#�(�C Tq�j�YSu*r.������K�<>5W179>G��gf^~�Xݹ��������.+Ը�.��� �	Y&Ic0mu�]��;LlV���ֆ]2a.�|�K�FE[o=�a4�X85�=�%�P����V/AK�Ndb$���
���(2�R��t�b������ޜ��R�~�kbs�ۦ�]�{��&S��Rk\B\c��#��o��x��cK�\ۖ�1̥܊ou��p�rZȠ�xu	焝��9ȟާ�F��|nG|Wo�bhp�Y��`��sb+����IK�h�=�6{Ǚ:_���������ߍ����B�"@sMGK:�`P�Q��Ls��A,p|��{'�ڤW�/D?EWp�c��؊�o9M��
��M�'�c�{y�z��e�#�F�l<�B��]O��%۰O%��<r�e5C�f_��!>�ν���g��_��/gL��f�#�EgN()-#\$�\�Y���DB>'d�f��d?���@4�7h�
ǉ9���x�5�������:V19q���WxQ $���%��56��	�2��ea$�E����Ғ	�tlRh��`	d-f�Ԓu���:&�h�S�3��я.˨��v�ٜ���j$cT��	�$7~U4��Βy���&��=���Y��!1b({�o��rz3Pǌ�:֦�<G4�R<E�e�̼螪oJ�e�=��{�ތG���#��Mx}I�����G���1[g���X��p��ѥ,ߋu�e�&N��<.Y�WNH�k�|c?��M�
�t>�,�s|�2#b��-j)�������o?�ǘ�}�U�ˉ�V.f^��q�`x�9��K�!m'�������7�-�QMs�E�`λ�_Nz3
?�;�e�͊��~�]T$r�Ɗ/U��
}B^���c�k���~���7�jF�.l�g��^pr�3��+q#��)������{�{�H��C���c�L鈈�B��\�c���ġ��q���jh���@d^�Ѯii{���;p��e}w9��l�����YT�'_!ߚ;���¥HfH�+�2k�5�ASF�j�ʙ·P:{���s��	��d	��pT��!i����x~p󂭡�RS�R\o�"V�XLq/	@�U`,0�������""����*܍u�P�xC�|A7K�e#,�b�m��:��*�8�NB�������X��[���J汁w?���h��09qװ��~�g�(�5�׭�F�J���_�J���b��5Ƹr����z:P^��kϹI��\��7��������%��|�SB�/�[Q��"��ƚrK��T��(�R��T#����-K3uwUi�4_I®g����x��t�S$/�������v�"'V��c���)ʮl�R�Fp�I�xrQ'f$��[������X�%Z)	��t7^�RƄ��g��:_�ޘ�K��������.���*�|�!���K��s�?��Rl9g����fr��F���f��J�CrVZ��_�S���!�Q�̛��D'~�A����W�E�pP!.QC~:�/�y��$�c��3��4��֋��ULM��W0Q�v#�C/�B�9��q�=�݄	 S���E���}�AX��a��*� WMa��ə�qOu���EDO��k�ء��NF"|V1r�>�R�ʨ+1�T��@	'��x-x��ˏ�g�ea�{&z��6=O5���p1c���X+���cQ9bǆ�����dj���[���d-*b|Hvցޫ��i�zeG	{i�*.�P�a*`��!���]}߷NM:V�hR��~�
�v$|�RP����(����'�c{!��8�[z��!p`�����B��۟�֚�-T7!��0 ���A�Ԑ��@�$�9	��#��AV��ZO�TL�����N���V��@�2�x�M`�w����@T�'��B|�T��)��J��o��))��9)ӢD��s�a�!8t��le�%?'B��p���?�F씿��������_6_=UbkN��Mj��Y�d�_|�{1D99k6��Z8AM��ƪ�����rF�Aq�� MWZ��m'FM����;-��<|��t�mN��a��O߰�O����O�',���;_�h��u���sm��$W�S�HĊ��ԅsv�wث
�� ��2E��4���a��y��ܖ���䒺���x���X�>/�X������w;Q��kG��J�ի�q �6ǰ=��I�u��F$���س]8���3�F�j��)�/!ݲr��Ք��4��l��hgf����c�&�IK��6�!�Q0���x=��]=���,��d� ������0;����=��i�@w����sk).�sOvA�y��W��oh��6#��Mbۍ	Fm�����F�F�2��PK   �X?Q� �h  �i  /   images/27231162-8669-47ad-b932-3d7f5563edbb.jpg��UXO��9	ܝ 	�$x��0X������'�Kp���,�2������=�=�ݷ�N���ߧ���~���6����hhh�/�.��
� �ٳ�ʿ��W0_`bb``bca=����������O�
���+BbRRR\r
2
"R��^����̗��/I�p�H�?��o �4@1:�!:!�� � @�D�� ��@{�/��X/^b�����
���Y�k��� �$b�yN���ɕ�?8���l}/��4�E��-�%69%�kV6�7o��ED��?|��WPTR������7 �[XZY��ڹ{xzy�||C��#"��c�SR��3~��,,*.)-+�������nmk���������/,.-C�`�;�{���W�k����� �h�G�?�"���:��Оy�ׁ���9���WWb&��$�I��/�4�fn��d,�[��I�e���R�
��tA��h�&� x�*�a�Wk%Q�Y�2�\J�7��W#1,�\M"M,��L�2�h���i
W���Hb�B��7�\����T9*_�9���P�?0��??d\���d��3��)M�j
�� �K"OT��/��"���q��ю@����ľ�c�bT��N�;�3-��݊�z������B����,W-F���	/W�&	�2�$��;o�<���⩐{J�x�|��llG&w���}=d�O�|��' ���Ʊ9�ҝVഁ���n��$"�Ҕ:�(�x%�%I�j�m�]�f���8Ng9���+	H1�BP�ޫ#�y�.�$�7�����F7��SK�EYB�+�d'%i�s��8D�=��=��I����V}2N^u[��I{�iK�_,]���W���u�M>l�
Z@`G����Z��P����> �	��|�V�[�b=6#Xb�Mj��PY���D�hD��;�}���|dEet�ox/+M��_��_L!=Q��I�[���I�IlOB~Q�g��=�g%�T���hN�o�4R��#O }h���֒�=u��{�������=�����f�\�h��ý�x02D>W;�J��rJ_ZN����S�oj����m����~;��R�>1�1g-#^��p�5��=�"ˣ��t,
cކ�h����"��ۦ��-����ͣ
ۄ�>��� ���lMUmӕ��C8�i߇ms��S�V-��_��y?ϝ���M���"��Y�%�P�d�X[�Q2e�����5-eC���~X6���bs.��*��>q���ޡ�"k�a��I����՟r���Ds]n��a�d�����D�t[��=��k�2�*��=ȗ�L=v㌛վ���j�P��ꇌ�g=�R�#�����n��>=��T�Ŀ:���tH��o�Wn��Y�}tvD=��<���-GV�YWV�	�
i�+�J�?������������N?Ҙ>��S'W	�9�e��D�[)��i�kҁ駡�?�;t��d�+��T��~����
,O ���;g��{t�?��Ϥ?���K��o4>6l�[ݛ̞	%F���uf�31��L�l����'F�c�<���_�+��^c"9�Ĵ)2��7��Gn�H���|+�x�n�c�W���<M\y����NW���KDzqs����|ܬ}*[����z�A+������W5t���3�{��{�ˎ-��ݟ'"�PCÊ��d||�/�w�u��˨~��G��3���_Z��h�)�$���k�����$����)u)������ް��n�����^uh(�4+��m
�~��cJ�P'�`ړo׿$�X�?��(����&x���a��\��z��H�b��N������I݇\�bҨ�-�}��D����͖o�:f��o�{Z����Y�.fT��ρ]�'7�� lR�	�}tI�ا��(|4� ��P�Z�X�����~8���bT�DC��I�d  \�sNm�-�ɿs1��Z�=��t��ߛ'v'f{q����ߣ��޿y�~%!�[?�/������͈j�7 �����h1��8b8B}�ǁ��wz _���];�!#k"��ȣ��ý��b[�^�/��q�|ӥ�����U���+�U��iklÑD9�s��7?=1�Vy��±+(��[߲3�w#^��+�������F�XA�J`���}I2�g@�}�&�ܶ/����.{�4}��)	�Q�P"�{[�	�Nx�V~;z�nY`��fS�a�ߡE6l�#��[�yk��)g����Y=�x����v�K�?\�Yd�񬤮���B^�����w˦�0I����dA-֤g(���81����b�E�?�ғ�H	�lA`�u�%-Al��9�?rjl�����#��6�jx�*vB|��<LC{l&^�Y���f�@~onE�+;!�z�ѷ��i��Q~����3����Q��z[�H
��v
T�-��"�������0�=�M��= ��"�9���0���l�����E��b�HqE_���#8��>�u��]C��ǜ��M����\����db]��I�#҆�9N���n��\�T/c��i_��v�b+�����[^�n�}�
"B�sJs���(�f��������F^�'�urlEBj)�Ys�������;h�=\7ԛl�w����y@�0�����"�zI�*���gD�ͽ�J����ORB���%z<�R�\��X[�1�'��uMv� �#���O	��/����~��<W�8�|,����R�`zo
�3���&��a�핮t���֗\/��5���~e5T��w��V�:�v�<B��%ٶ�=�u!��_��,~'/mO�]���~��i��s%J��cZRB�`g�k�B����������O�W'&�w\�|ӝ~�*��D���,,�u�wk�����'d�ՠ��]�W+鹏��`w��z�������Ɉ-ɟE���۔'1��v��W���.�84}�9m���v��y���D�=��1���{P��5�W;�����ח�߸��� �]7�={�{�h�R���d0�����ʭ�6�8AB��1{�z��J��i�+�!I6uRU%�����ʉZK�@r��3�sL�%���>�ܾr�(�ǉ�wt��VJ �
�iO��� ��I���k�6R��r��|�<��W���h[R��T$R2��������:��;�5Q�\Hzo�J�����;�:��n�h�+�[�7)]dE���4�]xjJ=�	��_c��],2D0��ٚ2@G�L^�w��i~KK�٩��"*��LE\���J���Np�h7�v��sdw��.��.S�Z-;��6�R��z���������y���*�o�χ�����~!�>�-�N��;d!%RbDo�qd1��E���C��������4U�Y�g��+Vr��s]���� K3��4�yNz��|,��V!gXpPۈ�&�_��8i����~���l��]�
yPw�!��3��}�Ǉ��%WlyE��Qb�]M6Ȋ�@��d�hP^jʛ�҆{�mG��0�[�
��C>������~��&�*5�2�Lv�W�גm���
!�O��>ښ`�K���%�(���8]x����'
�3�ǟc��F\9C+a��B���'?-����C.L�*T+T$ST^�_�԰��((	mYvRGǃ���E��xb��E�^:�r�q�I0i�Hm������Ii��p�%���`��q~���qH��h ��5����d��Kz�(�]V�KZh�(�)G5ӏ�:t�����̠J�0-�
��pL��3|4�S1s��a�}�g��QX.��2���I�c�<�S[Qm�T
��.�呇�\R�dG�Ĥw_��h��C�Ha��_���\�ڎ��t��}���-F�X�OP��=uzva�������u%}RM��@�!��� ����]��_�7,�?�sF�;"^ܻ�6n��Q�<���W�a��k�c��R�R�H	|�����Y�L���ՎaP��6x?%�.t��eJn�.<����	��X	3`jm	����*�:�Q�hp9���|#51Lqtv`��������H� +�:�=�9.{���>��g�$�P�w�`p��O��ݶ����b���j����NN�1�/RG�����kGW��RBPPc�id��$���Es��%6��}���Da�'a]q��qQұ��K��A��/��h� ��	!QNr)���H􅍀�5��)2Z �_���U�gU����=W@��>���@�n&H���N<�o�*{D����X�8�_ؚ&���H�9sV6)Y�3�Ni�b�pD�IO������ɤ�m�Qc��2}�\dɵ˟����z�b� \K�ub6��6����1C/�%u�͑�y��л�d��)���c�NJ�~$��Γ��WYh�ad��b��ϛ��~$Rn�A;�l��g�G�Ξ 6]�9��7K��o	�����A�yp�f��N�Dý�#vҵ�н�ս +�_ΏmhL슖u��ynOvp=5�������m�c���O���Qx[�Z���h�o��B~a
_��٤�p��Q�P�/��rSx�$�-�
��t��/�W�0�x����r*�Ni����aF�y��K�5��=�v�)��P�̩�_T;e�/�KDR����>	���W���Oݦ(�t�k�s��ɸ9"# �%�)C�l� �$Hu�sKuE���A�y7�bM��7���K.GǗ��03F��X�����A�7}��CѯЬV�ҏ!*��hsm�k��2��T�=��k�B��F_D���F�9Z�dz�E�l.�����$ٗ���Ae���!�*�%����6�o��hs���6;�%����7 �+��RT��ln�U�� P���x��$��`����P�\}�Ҧ0qtk_�2�ͩt'2ԎT���aͲ�FYj9��ׯ*Qb���uZn��y(fKe��r����m�J���"��t�����Z��n�� a�j��{ǽ@�C(wI�z@����XC�5��&>�󓤅�+�}[�/�D�5"~�Y��d	�v"w��QS��x(�$��@L�.ɂ��UE"���i�V�i��I5ez�㑢�|�=��G�8d��x!@��Mo+r�k4t��UF�kٺu�g
�<%�$�9��W��/w����H~�*���|��H����ҋ|�����F����~��.�˦��m7,������Z�D�����q�J��̙C#;i�r����l���f�q(s���� �r�.������%b�2Q^H�W l�\L�(m�7dQш隦.پ�;����>��2m�E�@��ኁ���>	c@���ݮ����1��CNz˟��^U�HQ�ӵ8�s�����p�3����SNU[�k�0a���e9h�u�<����q�fn�X�=Kw��A�[�{+)�k�q>������7j�M�.u רoƟQ�ܚ��[��1�K��Yq���:y���Km�H Al���E-����`�3 ��v��D#R*OlE[�%$�{�Qv�а��<q���cx2(c�����}�.r5~��D���v��x^�?�v	��W�G$(m�d��X��l��K�9��:����I��]w,xT��dn����I"2M���� ��F�K���Ȓ?D����)���h)����rU]wS�}}b������~���R��oŽ:��L��&U��Pk��a�1��J�K�#>�/�G��bP`媳�vNk7r-��v�L�"�K�mKV��!�6�l����#�nUݝ�d5�}���^��(�^��W-�9'��Gے�N��T�l8B90��H��	���yhࡺ�tq:���������/Z�Cs�k�{����1Q�O {�c�9�dNHz53�Xk���~�Y�Q�n�d#ێ��
���̞�x�m���pt�`KA�O��� �癇(�/����.޿q.�?$�CVY��W���K��-����vhZ��=k�aL'�W�.F�ي+�{6K�-pa�G�C�D�\9c��/T�h��J��$5`�*s����ܥ^{J,,����k�g��m�]�:6�~�6*ENis`�Y��Dd�w�0��r(�h`��$���Lh�Nqm1�'�ؿ4��NĶ:�%�t3���p%����c��O���Sz�<�Q04���6^��qԄ�u������9��lC-����Q���C��n�G�' !���i̅� ���u����ck�/�DX���E[r����ޕ@�EVN�s��\"��v-���k���.DX�T����	w�<&�y �-��P�Md#�ܟc+Q��PH�n�8�"Ӎ(�	&���9`�|[� �9_6���jutR�3o��L(!^t��嶍��y�x�q�hT@= ��2InI��|�	S�՜�88i;y��Nb����#|ɯ[y@H���f�J_{qµp�Im���c����>�b4�@�>Z`}�
��mu���pR�05߮��VU�Ld� Z*��AQ�n�k�j����¢!�2|� k� �z�����qV��*�ظ*C\������|	#��KR���ν�@�)Z�u�=xO �f�x��_��T�h�Nq?�ũ���|45����j�(窩����zl�Lh���S�9�
���G��0���A�&���A�<���d3�K6�i\q�ȔL�5�x4�iE��kZ�w��&\�;C�nxϠ*�@�t�����M��7�*�1��:DZ���v���,bFԉ�x2� Æ�)hA�7�4�[��B�r�5{�~��f���e�BjR��`�j��b�Vɼ��۹�����?z;����&_���.��9�b���stP���d��HW֚����AO,�&E�����˟ �l�A���(UI�D�"S<������Ԝ�"��?nQ�����e%&�>Z�3xMJm9�<д�!'�4ۉ87&��[�Mo�R��u��%e{ְ�f��`=r���q$� �R
�d|�|��ѻe���Y�\}���s)n����:\?��Ж�_��ɉ�� ��d��V�ǆ5>5�0�Ղ{��!�n�Y�Ht�T7ø����-�FS���+�\'�9� �-������{�+<k�>�����l��K*�~���t0�֔�rKi�Y�O
��e�a	N
�]~�?8��m�п��
`��/9�~�	�d<�2��KXu��!�p���i]=QB>�z5��R?��*⳼�؛�4�l��C�@�0�:'���2����	�Җt6 �e5�1�nOԄsѡ�>u~cd1�v�.1�	�h���/�P�ʧ(�2������r1|�˟^�vO�߻ �y���7�Xd0nO7?��s/��	�����)�^�uК�ݔSN����="�x��IVA�-�G�8f��~-$�~a�͏7���ѬG���g+\�� 4p����)� ��n6wh�le!��DO"�i}�2��#�R�M�GX��ϸ#�8��2��x��
Lȕ�0KO#��L��=<J���H:�)%`!�S�5Ԅ]c��_�ͪ>$��G��~k��>�R�X6&��q�:Z��;���sO�0t�ۺ��7pK��NT���	�7i��RX6�20���;�ͮ��O���+
O/�s-C�5�|(b,&˹4m��
����%��{Kd'+�9��~��\�B�yRa�"����� n���?F|�߼��@�I-�A�8ky�,�"��ӹ�40���x��Wbg�qQ��}�}Xd�ůSJ��w~|$�f�N�p$� ��Yv0�)�}C��k5Q���y�X.�y,c�Ԯ�/���}��{����# ��%R�j�>�l �HnKjmK���l���?0��߼��Aw�������8��h֏�o~�w$���U�h��P�}1�I�)J�����um֖?��т�qv2�$	h;�^Jq�ͬ>4��ʾH��\�^-}����v��L�#ǝ*mk̢��/罈������hˢ�o�?58��V��Q3)mw*�>��{�)i�/!wv��r5g�H:���n����+�P�����?�F����U�i-$b=W�3wY�u6��.F.�Ό��l.	��U���^��j�e���Ж]��6���5D���.蟏]
R����u��&X�
?AJ�Ȓ_�
\�^�^�L��.��֢��CU��.����Y�,%I�fN�}�%������5��`]�J�~���A��8wm����� /82��Z��ݐ���q�ϰ�L�o���(�
ǒ�O���/�~�g����R�}��Ƿ��uYYڔ�0��q���}�	��}[�Zp�DQ�1��7ղp��N+�0�4�&;�R���z%�~������M��9�5I�{���Y�9?�v��ۃ��Î������R��A�l���G޺�;:�^���i,�L�=�Uۑs�v�>�/���4û��I�US!�m�R'�y�i3��4�4��,� �1�ɗ���c�d�EUEڐ��H���v��C�t��k��,�U�ӏ_��>���>,[�xޜ�kv
<0nC�3Ÿ�p��v�|��b�4��,�S��d_�$�o��Fj�A�� �p�#����e@��q6��{����t0��ޯV�'=��#8Fr߽&��M4�_y���Ml��αe�����t�İ[$o�Y]�����!-~�5u���8�~'B��}�dEy�q�0aO3��D��Zi{޼�t���'A��˖&��5WW<�\�)L�=RK�m ԙOV�����&N�.�"����*�?�a�� M��Pw�6���rU��+4����`-��/,C�Ɍi+����6:���{de�l\J��	0�WO�� cM�Cy��L����t�"#�\�X>��e��-��؛R=�m�<6��|W�?���DR>@q��]4�#z>m->� �qs�D�ߒe����g	˻F��ť.�8Jj�Q����3��z��M#&/(.ȳ�ΉI�
���n���'��5 5��6[d�6��]��:]w�򙓳��1v�7}��M�A]Tۿ	�C!�>�n�h�2�>���g��Gh�L^}}�]=z�n*�S�lm�_r��,77펊ľYW2�y��V��@�k�B�'|2��4Dxė�m�i2\fݏYV��n�4场)����<(���.�i��<�T�#/u�ԏ��&�+]`d$S��/j����6����a�l#8E��>m:�P��o�Kז�Ӡ�X�8E
������ٴ�g�ƣl� ��z(R�z�h��M��F;���}��P�c� 
�}���#I��l��f`g�����yV�҇gA�c.�)��b�J�R9���c>�˖�1*��,��]�]z��9��]�@���u��'=Vu��)�DX��Aۅ1���$���$z�A�IG��їX'�[~θ��3�_H�S9#�F+�g,َ
f�Uhl)	i���	^(jD�H!&O3��>!g�{���턛}t!?d>�umT �i�����Pg,A�^��R�	����}��^�/��	��U]j�7����w�=e�hks��f��������=,� ۷+x�z<�E��-��^��o�׆J��OT�Oߋ=[^>T \
��v�/��|����NR���P�;��T���%[L���� ^���CDp%K���C�����I��m�[�:eE�ntՃ���	%��(�����j�S�E�M�}W��q�������1`b('��d'���0��+'6��I0>��9��s�E�:�����x�S���Z�M�y#|褙ؿi��M��w�)\�?o�z��B3���79�f��c_f�.����O��G�V�Y��E�vB�Ѿ�	 �Y+$P->ΧND�/����4Ց���@��coG��;n��n���+PȦ
o̞��Y���AM˦��P���K��AH}��ҿۗy�h(��5�
�z])c�W�'�Z���G�gb�b/�qݜ�t�?�o����r!�\\U���6�#�t�Dʡ,.=��4�VL4�;�;�ƆZ<�Z�s�5P�8X�q��tiW�P9z?�� 5 �͐��NE����5��lC?�ZxQ<\`��)���W��׊�@�K�Q���k�"��߄PW��r$�pQY��pyMɡ��k4swÝF�Co.(Y�O�'&l�G2�����4sK��C��1�����d^�%�~��]P���x�f��f1�����R�P���P����k����[8 O%��̈మ�����l�c2��D,����*�Zh*�4��"���c�J�Qm��NƷ�H-�	T��b��;���yN��c$W;�'rY&��Q������5_JS���bv�H"wd������u�����.m�U�#  ��I���:,��X+�AŁ��3+�_���1�\�� }��OJ�X�e�顄��)���������r{�C�`��7Q[��5'��5
O+� /|���X����P�a���fjJ���s��X1m�N��w�cf45���z��(ؔ�@��7�0��V�f�X�Ĝ��CI_Y��Ij�k��I�L��.��Y�J�ˇd��9���g��d�xE��(0{vO��f�<N5B�;��£Y�oj��͵[��J�e�Z)O4�s�t�2�S_��W?.����e�R6�`�9�PpMt��^��)I����E.�G�:�t�+8�����<ްY����Ļ�F��YPħ�V�\������gl��~�5C�l�CB۰����8<]�%A�֦cn�Sџ/���^�X�$��^��5�ͯj�|�tbƬ��h]i���c�2���cU��u���wj���e.u=��,l��ajSi�>�D��4U`<������j4����}+����M7��$H��qPP�^�1�K{Z��r��U���S���H��KZtƉpQpg����;i��Td?��xP�`y��I}��A��p�%�W7���5e����FK(d�C�'���P�C�|���o?z�c�-��p5���J�6}$�-d��^���x|PGp%Hʔ�M>2R�$W٭{���`ԉ�\�ބ#8�}��{Ȍ@*��|�\��}P�J%{g,��}��"�$�vO&'�+����20 �r2�=a|�y��μK?c9����G���;����/�KQ[[U� �;�
)(�'��	��9��f�Y���`Q�T�=�!��X�ue����r8�����g;>ã��b�!������O K�h�Tk��;s��ڃҩ��]�2��gǇ�Dt����W8(����_�iVȶie
$��UQ�7>$�,`�B��̯n&]�1ž/�/�I@�Ӊx�b��������3���2�)��?���A�-��xt,�簿�Ɏ2+��*okvG���Q��ؘ`��� t���4���уuB9ʤH�.��P�+A)�]g���<yD��
! ^���{S�G�}���4��p�.$A�^�F�(�%�׿��y6�Ҝso�{��Ȓ������\�.֦ �N8=j��̚��5@\�6FҨ,{hK%�"f�4v�8�5��&�"C�JC'
x.�s��!��c{����M��¿���Y�ug�똗׆k&.�ߚ1r�BNg��N)v:�f�Ν��`�]��̹�L��P*QwO�8���+;ra�ݶfu�C`�0~@��+k���P-p�ܨ�H�r����I,��#�N�q��Dh��y��uW� Ы��2]sʔ�ĵ���M��|�T�Ð��|�!�l h�ꑑ9Nl�T�^zp�{�J��A�#�u�>��$�U�f���.�8Xn���/�� A�N��0�x��e�{&���	�07x9Ǣ{1+�o�e6(�j-���0�Tl����@��Y[�w��%�<��v�^��%��e�'�U��v�t-��I� �@�
�%�9}�w�I[�&0:u;Y�oː�y�u�R�sByⰏ-]�������1"[�b��ѝO�a�h5�f�ʹ�uu��O��ZWo$u"���
*Gpli�P�]�quMI��xO�<K����5�U�y����2;3���8� ���wZD�(�PT��9�% ?,3ٶ���m~��Ƕ�' �X:���G=5Z����I����������m�ҠA%[[�� V�w������#�|mr�tJ�Q��J~���Nh����pk��`lh�Eƞ=�#�m��+�J��\�(K��i��
���V˄���^�����gKSާ/h��pP.H���O��d`i������06;�����
LW���;7:��i
�p�A�;�(�|V����X{"�?�~�Bf
r9$IM��S�g�?s2�U\��`Z��F�����s�9�^�G�}v�~��}�2�#Z��&JE~Qa��ӈu^i�f0�Sc5-����̪�V��|�Oz�Fc�ϑ������3�.c��Xsq4*���0	��o��_B����.��O^s�B?R�#8���@��#;a�?��9�l�����k��Oyv��K�2ۛ�t�0t�0*��Q�����;�;&|4�Sod��Մ�ۿ��B����3���4ו���*z��$�ݤlr�/��s0�8��Њ̗�<.���5���K7|�kQO7�?���$����
u�Z���M��(�oK}�?j��S#�w������Q�^��Bc�������ӕ����xd1�W��@Q)��A1��}�n��1���[���tҷ�"�(�G���Hu|q�@�T�=߬�TJ�|B�z�/<��A��䯧���@����8)Bq�+�%�]�p��r]3�[�S��Kob^l��)�igi��2�&֩����Z.GIX��'���ޑg�.bڑ+�ӳY��^}/��# ��2���m�,��Y1C�bC��]�sO �nj�{�z9�O3����e���T{'���r���ُ�E>(���z�٢�:�b�	6 T� ��W��i×����ƭ���@Q��K���1ND�L%`�/ne�ÅM�� ��-�����e��).[���yEA����Ӡ,�͇pE���f�ƍ�)j����"ٯ��֚�Y����T8����܊��������)y�eJ`���Լ�������?��m{/�̃��m��4�&�qF8}_����xm�ުg���W�[P��?A�M��EO�w�|6��0j˔����]��"i��N̥���߇i3%K"J�� /KK�L�O��u��}�6o�Hg}s��� �KxI�Chb	��4��}��c�Q�a0A>�­�P~ɇ�}*��������N� 2���eGp5��d-dU�v�0�=+~�ԇ���՟�1X3�_ZY1�r�|����L��=�Ǚ.����@fԝ�Hb 1�y��>n�b��t�h�T��֞�G�b��}��%K�����Jr��L@��4�\8���{���c{ʇ��b�F�=U=CϻzM��f�Z����|͗�]���XU�<C���?�3[VdO W��og�F
~�ދ8E�J�c���˂��{����^U��о$��������,�RΨ"6ocV/v�P��ˇ!��H�{�Ĺ�w!��P�V(y����������R]��b���Ox��u��|��+
�M���g.�_�D�1������QGxr��(�%GDf�
�T=N���ōXX��u��P5�z0_��h��;�1i^bԧZ�as1%�2/�Rc�e��LQ�榵��36i��N��A����|أ@}���7T�� �O��;T��j84\3����`~��rc�9S�[y���6���8t�]h@�t�6R7T���]�y�ʤ�ƽ��v@�*]�4��*�}(Qh��4��W��ҥ�ֈ�Hgaga ��f��=�O��ݵ�W*�Y�><���A'�N���y�-Ͷ0�h]蛽٫���A��g��;v�*�����o�Q���iӵ0מ �AML�9�\�N7�¦���T
�Ad8]"2��!��*�ё�`
�i�n�ԉ!�3xYr������F���ΠE�9⊰h�]�u�߽��l���O��:�Ō��^��4k�F]�����w��杽mm�~虧_z2�p�u�.��}�xݰ#Hj�jʣ��me�Z�fv�����D���C^����Or�,��,]<ic�3�L�I�{���O�����&��߳�i��,�3�y��^���-k��dʈ�̿��T�%(�Na/�������P��Ğ�*&p�U�^nӒ�A���٨ݹ����kˋd
�"D;2��8�(�_���F`榱Ky ���ה���s�D��d*<'ŮwV\�����y����)A��n�D��ԕ��8<�I�Y.1��㘕�>�Zm���䀱F��t�;b"soÀ�a��%����8_9��?���V;8�S��l�����4:5�3����������q>޺.���:�R�跚~���u��+�{�¿���0�رy�	V.�Ùǽu�zU燔N��i��ה5�X�^Z;�S���-;�6�WVT_w�����h����5�Թ���:��UԪM;W]-%�U����)�^Z����&��JqI�2:a,%�����M`�^?'Oxg�"?�l���;1��U���l9�F����s��V���4�O_�Ĭ:r�b65|Կ����T��lW�$��|zD��-�E_et$En�/�[�(��3�Ky�`�'��nRax	�L�MI{Na\/2%YFd)�0��b���Y%ڣ�@�� �� Y�q��O�����p|�u�#7�]����XM��>���X���G�o�6n}M<93m���{�5���c����tȀ�Q4����d�c����<2<�UxU�}��25�����d�)6M���a�����K���[�R��y�
�)�\���K�w��x\=���s�?Ֆ1>I� /��㻋�2V�~�Fc���#P�|�9���{�6�����矮��B�ȑy������Ё���A_/��Q�/�ٻ"�]������r�zxf�T���[9�Mq���m�{�w>#{��I^"�Z��z����,�e����1g��p"�6d�A�����a�\�?I���������T��u�1Ī�&+M 8���]�������.����V/�EL�K�v�И��uJNDc��b-.O�N�hd�[��#ԫA�eVA��uS��TK�����e���z�Uݑ�i22���>e2u2c%K��/Y�\L�D,�L���ŧ�[z���h����q���$Z�_�~職b�=L�i��|��Jw�m�L���S��{3V�'��jm��4W����a�,.�q'��˥�j��3��J���P;�Gz��Ìd��!p�(J	7rR�G�e��dx�@�cZ���͝�L��T���`V�v�rWݬ��t5��3�Q�����c��ɍ�wM�ޚ�-+�@�H���� ��)w�Zs����O3��ӎL�N���ˎv1bf�Za�LG�K���<�{�b���P�����r/�I����8Bzc�p%̖?'P������Z��C�>0��t����ye����c���^��a?����������]xk�W���70E��ɟ#�!�I���XCBi�,���7�BvaV?�-�!;G*�!��H�8J]i�J��}t��jp�J{�V��V4�V��W�2c;(��hӰj���x���!�<�t��&�c9M�k[@1�o?TP�	`-�z�IREPxq��װ ��P�@����-E�הk�~XW������[�?��u��nM�O�e��2?;s�h�������g<-�ES�FV�ҽ�A�����8v��A}��f���fW�p3a5JQ{ui?��u�ZSS�~��ڡC�e���#�^)�[��^�v}-U&H�i\:���L�D*�d�g�cڵ����xխ+me���֛8�u��cN���g��2��-l��� w�>�h�g����y�ȓ�2�=օ�ef��_�h��4;�^_���I�(O����B&�҉�!_~;�5c:�a�1s����TUu�5��9�O�;�,��"�ZI�N��ʾ2��P$�>\��u����@o{�c�ǟd�k��%��Nz����78Ո:ӫY�3��m2��x�gM�ے���&��|f�:;/��ƿ�U:��l�?+j5��ʫ�M/�)l2?%�O�c�(�n��c��]�+J-�@ڹ!<����D�is�U����)}�KDs�mE�#A-��1��y���R�Bz�CեG6�k�y����ڳ@��^���yܼ��^�VC7�J�����ZkOC��̕�$��Lb���?�����J-FJa�3�k1Q�+?(�׃P������1��B�5�YM��A-����6v�y�����V�A���n4]�E�8��t�w���Z���YV9$he%f<��.�hT��K���.Ɨ�0�uH/�(,�Yd�4���G�-
�q�.6��|b����`�ĭ��j�5�d�%�,�4̬�2��Ct�I0R%���i>3�u�E�tD�p9P�ӡ^�N�r�~a�23���r. ��F�w'�4��m_;�5��)�F�D`G ���>�^C�n��呢�gv9��j쪽�$��q�����`��N��j�'R{��X,�f�F�h�?�&ݻ��`g�B��������[��L�ѻ�{zQX����Z��ml`���A}����23j�9o?e��i��/,o��U��̊U�<�,̭�,A#�K��S��A�4���58d��hT�38O72m�y�?���v>0�c�ï�Koww.����g��帖%F�A �X��G͞+��������n4�;�r��m%�����v夸���셕ry,'�.��B�qS_[k0�$��ͬ�:O���|�!{F�CT�E��H�OJ�i�C����]�,Q�5��#h�PO"�>b�´�`54�>����I��/�r�wZ�;�I>���¾�`7ez/��Vw1܋��],�0�Oޤm�yE*��n���8܈v�*��ˉ�z��(�՛P��ѬE}�(��Ӭ4�@i�]������/����2�7%��ɗZ��Mb�%���&���Rq�K���ญ���2�dbcV�k������Z��v�Z(uk�J����6�^�	�T��<�]st� S��� ���V{蚝��U�淧�umR�;�`<[˦+�� A��jY�#�&��ޡ,������mNU��ye��Ha��.���+�;S)qD6�~�[K�ؼ2?�R������D[�-o�ŕ��a9Y>bZ�j�W])�_E{�@�O_hsk��do%ͽ����*��yd,����!�Z8d�-���� �n��;��m:�($I#���[�6FI*y�Cw`W�O��#צ��� n��5�P��������BN��l���h��sH0�e���a�5MCM��^�.u���H���I�\-sQo+k:#�sM-�K���GnXn���&}R8�-����^�_��u˘�H�o�3Xu	vRB��ܓ5x������;Ȯ�-���V]!onf����w�|=$r�y\+<А�%�����Go���J��|io+6�I����du�X����\�����m�c�e̶�v�Z�/���ĵ������a|�o�N��S����K=�G�C�k��1;M&�7���nb��_�WKԬ���f��,�Z�4�}�R���3�m�,�U�/.�i&��W���n��5֗�[j�z]�0*ˤj�o{	x�E!!�K�;�>�X쌞�u�ͽ�߄�K�Z3�WL�Y,�L�\&B6s4l��1db�-jV��Z��\ڋ���:��ꖋl�F���I�]�VD�����LrT�ou#�ac{'��R[��?M�E[MN �.����Y��*Ĩ��BT[�H#�5Y�94�n��h���kK{ˏ^�y ��u��U2�ܪ�2�Kxդ/ÀK�Z�[�f�� ��%�ћ�a�N�K�1�f��SG����1G�2 U!33D\=ik�\]@��Ŝ>':pՃk1_Y�n~k�_�5Y<�,��B�2�%$J*i�[i:��(�+�PR�J�%���y��7����s)��wmX���c���[���7��q�16��ƞ%�-E�k7�.�k�yd���< ��Ii��*��"����T�����Z�!�{..#:�������0�|�v�h����q�s���ޱ+[�}�m�-緕�y|����sq�bĸ`�#s�F�A��mn�'��L3hV���Q=�V���Z���I��֍fGQ��_T��ա���M?M���K��a)c��֣th ��T�`� �L�����I>4Y����Γ��Vܭ�����0ߩ���������1�K����b�.����J��O�b����),��	v��*�J��)$�X��������kq5��vSjګ\�$�ח� �E!�a�+t��Lp^6�<s���?�i�^]�5�o|gvB4��h���[��� �݉0.�u8��*6ճ�oX�x�_���n����4C����Þ'���x[T������$�7n�������Ԗ���]�w�v��'��/g}s&����� B���O��ao��m�'����K��c#Ew}.�.�^��M�Iڪ��|���1�� �o�����? ߖ}7Ś���
�E؏��T�g�Z�?�x����u/Ͷ���Y�X|���D]�w UX��8W�����L��b"�������>,Դ)��L��<?ذ�71o[I?y�߁�Z9�L9�6�5W�~&� ���]/]HF�yp�]�:~�w�g����b���w�55��W�ŭX�luy�=kV��5��3��󳇍�����+���Flu\�%��󭷉4����p�q�q
]�x������qckH�^-��=I�+�'I�X�h���^ũyV�щ ������?1dU��'�6-r	4q�o�ӯu�x��z�M��R]U�kx�IH�ڢ�*�)Ǜ�4���W�ϴ��Amo��b���i$d�)��<`z���=�����9sg$�c6����z���I$HZ&�B&�eQYX��T�-��N�Z>�n�[^�� c�iP��0��!�����H�g��(���6��b5�%�ֳqmj.�o���oc�5(����6,�ǧ߄!Z4�2�|�`�ui4��t� ��E���i����薖��K��eeuu{ď�E���h����+|P��c4z������i ��U����$3G�2I��P	U�x�$�����9�k���W3G���id�uucwዧ�1��y�KVGnAN��-������|ꚽ����ý����������09����$�Mf�0A;�gG���o�ԭg�M���:v��������^��O�B�� �U�ړ
��͗�.V�.τ5=JI,�����v�MJ����"kP�%��v�U,�c*������Nh�����+��5=>/���K9������Vx���e	n�r�I�!�Oi��ַ�,���n��N�cp��f{[Ԇ��tA72�{�b唥]�Kkح/�HE��^^�q�ͣ��S_�1@��Z<������:e��$�wS����6R�B{}]<���]�=N71��Z��B�eӒ�&��&���w�,���Ӗ�QK��K5K?Q�/7��ѵ0.�.|�,{«p�n��o.�;	͔�,wvO�(�P�O$4�I�H�so<���蘴m^8S����[���2A�MH��Zk�ed���2��F_C�4�
̿�����a���H�����5�:�ha���B�q�i�N���"�k!e.��e��X�Zhqˤ���S�ѡ�hon���7V�i��[��H@�q��e&�XGm�ɘ��L]R��H�;K}Slᮠo2��Y��Hq�Z��y{��Vs�bO�G��Χ�ɹ?���m�ˑ�Y�䋶��&���5ϭ��/���O�t�s����̫r�j�mrAM�u<Cy��X�*�	���b���-|�R��Omqn!�Y��[]�� ��؍�6��v~��{3a�Mf��m���#�.�\n�u�X	ss+�k�A�L�ݳ]EҴ=&�Z�/J�\�]Io�=��?v�xg8UT_�ݰ9�zOxV�P�|GV7��K�A�d{yP8��� 7H�I.�7Jm�)�nu^1�&�s�0�z��t�~6�V�Y��J�q.'��Sʯ�������I�կ�}�+o:4���ºt�#H�oE5��~IVO*0���MW���Ss㏌��c&�g�%��K������Rp���2�X�s������ ii��_��O��ºt��jM�ۋ�8 �g%W |��]8J��8��;B��o����c�BjN�%���e���!|�4�ߨ2c�W�$ծ<Y��:���Qԧ{��$��c�>���T0�T\uG�Kv�='����ߊڞ��N�����%խ��I	R=����~�|��e�c�Γ�KKg�N� {-SO�0ZU�'��p�_�OZ����o�ǚ�m���L�\�5g����:�,�+�x�/�o[�,�/�&�H�:����@
��Q]��^�*r���_�ŕ�ӌ�����3�[�j|y� ���Y��vA�y1��A���� �CLp���6�?�χzU����HmD���F������؊r1�܈�~d���h��h��|�ci+ t�nY	_��Gu<[J$}��#��oݳ�>,�4�+�=�='ŖWok�IiӼ�Ad��)�VT' �3�T�ލY��b�%x���|C��(��>#���G�Y�o�6�z�G�6��c1`*�9�A�i�c�����'��$�l��3�ܒ *�Fq�H⟭x&�߇���kj��z{�2�%V����B�N���n�.�ݕ�u/
ދ?������,* :&�#UX$l�.d$.!m��ߡG-�/ ۭ����ݣ�����D+�hfk�Y~�;��UK����O3��H�jf�-a������c�⺓{�h~�w8kX�Q�|߾�6��m�͑Ğs[#m!�,~v$i26��A���Nk��/Ï6�����\[�¶&i�C�;w�W����o;X��^I6`x�՛��������*�Ig�K�Zj�<�C�]�o*�����6�ڰ�6�s��Kw�_�xi����S�W��K����Ye3YĖ�H���*���Yt��?r���E��o|R;�0��)Zi�gH�HRTH��1��ޮ���6��]��m�Ė8�:kKy��i�����.� f/���f4Xh�e�����g�ٍ'�^!S��Ksm�V�T��� =?r���tŞL.�7Hj��<�Z�u���5�BdG��;�e)}RՄe�y���3�ce�q��uX�����k�O�5�l��>��S���Qk��yP���Je����f�>�k� �PAv�nB=��Fe��m%���f�������I�-Ɲ�_;k6���-��7,��SP�p.m�"`���fZH�t�k�\�}�����
5}2}RԼ�H�,�6bx#"�c���-2䭓6�Y'{�w��V����3��-%�-�� ��������XgD������F��~�$wi�x�M�hf�M���I#ki�2�x�=n���&y͏���F�A�i��t�紵�dXWȷ�1>��,�����y�6�P�|p�Iq1�t�I����O*�"���3�����p6��ЩZ�g��/��8��K�X�^	n����?�(�!�M!Tā������� ���w�x�M���a1����� ҄j���2V�1S��r��$�=j��.�k}g�7��dk�9�����d8��2'��EV6��϶w@U���Ş�/��gL�S���c�Ffe77R^V��W�;�2�[�����g�<U�kZ"N���ɨ�N�f���R0w*�P�8ڀ.�V�Mվ/�Uxu-��/-#��t�;�	���}�
�nY�����ȡ�e���ƖI]��������Z]oX{�/􋛛{z�%��3���8�̲�6���s���P/���Ҿh��wz��x����'�cq���|�����Û�^�e�����ڕ���3Eo�n]�q'5�}s�j>"�/uMZ�K�R�S=�̇-$����J���%:�X��G�f��rD�qݘ���4U��3#�c�~tW�U)�v|tqL�ό���@׋��\�1��\B�v���8#��k�>6D#����>��eT���=���3�k��S����<�I���v}{�#��	5����j��W�[���	a���}�#��g� ׺���:^�"��S�V����H�}��T��2y�|�i��y
�X�Vh� 1gYP1�� �`��'�+�ٯ���?�<%�R����4o.��?,i���Ì�A�~}��m�������Vb��uv=�!��:u� ��y}�\i��[��M䵫�G�H�EA�P�.6�R�	�,��I�N��}�?l�4� ��n�͊$ze҇1����}���KбV`������ݴ�p[h����	4�y&f��9�d\��j�bm�m�
�9�sE�7�~x�h����N�ZK����&�m,���L ��\��g%(���>�N2�,�	>�����7���RG(�osw��)��o�kV$��-�#&y����L�t�xoU���I$	w�i�v�,�s�D�UD�B[hɯO�:U�o~��Y��g���ؙtˇ��U��Rb�M���If8b����w��9��~
�yaȗT�.�'L� y�.r!=�6���OZ�aܽ��i����H��o���[�:A4,%a<o,�ԁ� :�T0��j׆�y���ܾ`����e��� �H�$0%L�Y+�ǿ��5˕� ��H�u�������m��P�<���C:��H�pG�}ῇ�#���9�5EKh��\�b��*,�*��<*��K�(G໤�"{湖Gi$�dX�M�^p�)3��,e\�ۗy
el����C���\b0������H�!����+r������Gז6]� �l-���K�9���0U#�����:Eլ�.��a*���]sv��4orT�X�v� &�$־ x�7��j����#C��=��4Imwem��H�[o�s.pd��^YK�-?	i	!ߩ���i.ojm0X#��aQ�YT�ܒ��i� ~|>���JH��o-����u�<�X�m$��H�NsXڗ�jv��n���M,�.5��<1i<�_-1�Kr2*������^�<]��rmCœD�^��B���Z;Kx���-Ŏ"U �&F�'�~(|D����r,���m���}2-%��$��f\n eTß��+�gK���կ�S��@�Ơ�!�]đN_ 19	�1�u�_���w��C�����mR]�� !<��,��$k
"�H	������yï��⦫e�hI5����\XT�'.�HG��Cʻ�n+��'>��|�^�jrC�ٓ����u1$� gi��Ir�d��<�,Y�?�|�<��o<?��D�-O��C�FO�@kn} C�G˒+������w㟉��u���n�g�4kb#���j ��� >�,ɥ���E��b��C�2|Z��:�ٵ�R$���>Ϧ�v�X,m�ݍ =q�ǹ�V�g�\������rF��dV?�l��(o�'�x���J4�Cc�f"�Gy��h��(��h.��2:�A��x���Z��
u�ʵ:ߌ���?�]��n>��_������y�2� \MMS�˦�E�[S�cVfm���%�
���������t[�m��xa�W�ڤ��֟���b��h���*�aO�W��=��s_��հ�z8z:^*��eX
x��jT�/c�'ğ���n��7?5�kU_����o5�c��^ ��`W�?�	\xGB�Ě�ƽ�h�E���B-CI��X����zJ>Oj��?>T�����?h���Uǌ��b��"��W��ۢ��PN��f�I@`{s_��q4*�)6���V�Д*���?�� ���ٶ�q>,��)s�\o�)��Il�g�:g����?~/x+�4v�>�-5�+l��?K$7�L�XjC2.d+ 8�@?9�l^�����Hֲ�n���1_�qQ��+F��$O1�lA��ʟ��+�\NG��)ƪV�G��̪a[�g���z/���H�֮�'s����E�������e���˶�3��?|������QG�>��[[��g��"�aWF��M�)=�y����Oû_��(<]����"Ss�c
�޼v$��^����C������H�O�-A���z�M����j��F=c$ +�1\1��/u]EG7�5i||]q'�����Ko�)���H���	X�P $��8��k^��Rms�w�B� 7PyV����F|���^����~8���(xĪ�c��o�.?�^/)O�eh?���F�C��:«�Rk~kB���o��'q���y=kÖ_�����^8�2WL�n1�۫W�_-����̷J	E�# X9<Etm�x+��L����Xn&�y"�f�OtV��E}�?
i� 2�>�1�%���G � i|��w�&����<�%��#�� #��ߪȝ ��� ���G�+�E_��-��:O�Ox�T����7��P��Ŧ���A FK"1 �
�ҧ�J�t߃>�ї]���Xx���ɩx��(��fUYbP�Օ@�������t>)��<���u�Ž_Su�?�qX@J� ���:c*���i�_������M�1�?�I�jdg��F,Ԑ+ӣ��+5�us*4֌�OM��%n�(����L�+N�(���'F��3$vDy�~f�;��s^%������"��ox��F[�P,zv�9\�Z�ڃ�!��O.����/x�ⶮ���u��v�I1��*,�H�
��k���y�+��RO�_i��Nҙ��͹����>$x��5+˭{�:��i�$��X��1�~� J�7���-�kH��ºo�/\���7%�r�[�R��,A���'��{~�i������
�������]�Y��1�Pơ4UP0 ��g���}Z���ۖӎ"��?3��%]x7Oy�e�C��ɛP�cIch��� vW#�Ҽ�����4��/T�+_��ѵ�#)!�q-���3Fxa��~�K\F�H��pU��{W��y���>����B!��R���:%<A<�X��e�2;���Ǔ����Eɴ�Y���Vh�6�Ym�cBB��Iy��S��h�ثBN�g�t��G���(��}��5ؓ|�e���C�B#����4����u��g���d���v���Ư�V򷏵) gm��#�y����k�#���o�s�֡$�r��б'$���_'�dr��T+a���=<m�UTZ6� 3����^k��&��l��{�ԍߔ�Џ0�� r��� I�֣� ��6��{}.���k\'kc�k��a��_ǭ���ԡ�e�Kv1��d�� ��s�¾S	����J��>���%S�g����gƚ��w,Sݬ�;�y�@VB]y�m �@ ���XQ�~��5�֧�]_��%����su4ĳM+�gv=٘�OS�yѝS �������Ҍ$�J��b1P�ۉ��ʻ@⡒ܷ'ԀO�ֶ�K�7�>�Jci�����j�.�*���Z��E~�8�긱E�����y4�s�/��*?�`���f�凋�t�U��:lQ����*)�8�+`��@�U�� e!�"�݅=t-�>`��d��W�-��\gsc��*x�u\t�*�������]pdS[B�De,Rfڱ��ԿeU!�sZ����ߨ��h�ԝ�9�f�#��X����o�->x����t��\���k�9d��RFY\�~�~����i�,��M&�+��а`Aο!�H�0)�t'�_ýz��8�[�xgė����w�?C_���LuO�P���e��0q�R�h���h��yeu�4��m� �Oa_�� ��ǭ���ׅ�=p�{$_�^D�L�B)�2I����!�;��X��*�{&����}@�+�Ok����<����7'�j��*ة+#l�>X�N�(���t�Yd��n�V��.��,�h����E}�j��F���-N��V��}m�|(𶹬�q{����I�3��2N�9=�u�>�H���*	� M��� ��Q_��R4)�On�V�Y�(��� �>�
���=on?��t������l��=��� ���Z�����*|�
��˯�[�tn�|/�@ơu� �kP���G&��� q� ��r�+��U����J����g�1ے<6��{���ԮzO���(��j�d�� ��QYʵ_�y�J�;�+�"���T���8� Z浏���y�m$�)��(���Z��?���T� �}�)�xsH�;t�� n���6���4�03� >��QY�j����T�� *��鼛RDV6�B��j��C��,?��� E�V�U����T�� *��<�U٭2@�k� �iD�e���"P?�W�,M�{:)Ѥޱ_qb8� -?�V|�UUzQEsT�W�����aK��_r4!��Xв���W��mF������h���"�������4�U���b��z|�ox�,Oi�&��+�թ���Th��^�����PK   ��X&�n�-u  #u  /   images/2a76cb7e-09fe-4529-8dba-ea35a2db28d0.png @㿉PNG

   IHDR   ^   �   [�7@   	pHYs  �  ��+  t�IDATx��i�eו��>���5qI�)�����Zjɲ�n�q�vv0`�F�8@~�W �� ��@ ���;Bl�c��lY�Vkh��5Q�X��*���;�ag}�Z��[Ū"�������ޫ{�=w��^��.�w�ߑ�w	�;t�.����%���������?!��܋?!���������f)�K�ҍX��$�f��aW��ti��������eZ��h��m�Pѥā���4�>B�"F�;��	]=���w$M�y-�16�w~O�����}3d'!�<}_RJ�!P��شꤿ�,;麮�$���^�R����x��<��/,�!�o��cS�s,�3Yv"��p���������g�ﵾW��]��|������ZF(�;���_�����voؼ��'����<��^�xS�����:����m=oT��zۮW15���?��O�/��G>��{��]��R
��|��yp4�ԬGd����Lp�LP^J�U����2OJ�j�Z���ܕw[���%N)�a�M�OU��wR����r��V�=�q7���^`c�B�u�-�e���E�UK�1�N��t<AY������?O��Pw�L��Z7��J��?��O������؇_xO��fJ;%�?�u{>���R<�*)�[�U##]�|�}Aɪ�X�:�(��0�T)�-u���H+e�FbYIݶRT����\T�^պQ��+{�R�s��N��b�ڵ��Yא*$�õ�_(*}n��f�w'c}n��Z*�M��4:�AQr���
����\��(d�X�`�=��jy,{{{�&�S��hC{n2B��~�?�߽��?�_��?�G����p��C�"�\K��_�ڏ|�K_=�T�*�p��AEj/�+I:��I�Q+�+p��WNQ:�J�g��@�Sq�;#�Z	�7X^u��!'eҶQ^�h*X��ަ�k���X�F�&���Iǅq��V��D��e�L�s]Le�(z�é��W���!sp�A����p���\�ZuG#PM�Q�BJ���d������?����������,���#O<��E���	�yp-�X�p���7.�&��+�I�9a���:���N��AcO��rp����:ڲ�{��X�zS_����u�S�G�h�D��c��C��(%�M?��.�%D5�s*��.�b��F|�J�Y��5�˅
���u�A��U����ua�������Q��T��
�`��*���K]���MƲ:�*�=p]�̟솃Nvv�<�ȩ��'��?��&��7>�{���b�����B����I3:�*�����R'�ꕜ��WK��3��Vܢx�:��`:�W`{��K�!J	Q�x6;��Ɉܵ�I��j0U10 �g3��N�}��J��8�b����#ٛ��m���RU�p2���U�RNw%NZS�JP<{X��jiu7�tqֺ+[}/��H�[��ѱ�t\A����9���nԅ�rWE���jmI�dн��ލ��L�3���^�*G?5��;ҝ:k�Qֺ5�:���j�(�Z�b�b���\��3O��~�S2���� 0�=��o�/��W�{Z�������z���S�ě�|����}�'����:�����ȯ|�k�Ra��	/���mQ	�ЫBŇ.�O~��ȃ��r��8���ي�������k�+�(
׺��x�VE�B��خ���;������s��1Tqb&2����/��\x�2��L��X��Qؑ3e��꼹ңU����]�U�����ʟ�����^�x�g��S����V�\�h�������d����}��?%�#�M`��u�S��_��Wd�� k�����X�܊�tUt���'��B���u��y��|�+kG�~_iַ��P/����b-���yLfǍ�'%mݵ>��?'����@5AJ8%R�J8$]U������O<+O?y�*��~��L䗿���Z��SR��c�FE��.��\߇���E�Ͱ���庫�������O�����:Գ&TS�I-�N��T�$��:�� r��z���P&�\�*U�+ǫҫ��Q٨� �����o���"��\v����oQeլaK���ve�JXp5c9V�^�J[wʸR����������7���Te��nqM�����d1pfT�^E+�F}��;R�N��j��@��x_v���7��u)'���t��C[�h�{B�{��[h<(�wKx\��qX�붛�؍nǵn�b�#�N@_P�<�a�����;
:%Z�_(Q[K�����Jf�R�Q��@	�O,�B]��M��B?�&���ٿ��U>)g���E�2����u����Qί��׋����ִ<u�J����	S�J^	Y@q�+Uؓ*ȴ4�Qk��t��2֕��XԎU�V�5�7�_��M�����9�,��0��r�ݍ���jtn*;<����6��t]] �vQ9x12W.�|��jjI������T�UcYB'胋rQ�x*W����ZjԮ�ܬu⥚���tc}�~��ʽ*�'J�5LX��P~귫�[r���V*~�c] ��n�1��8W�%�܎>�*S�C�;X�:�k`�" "�`��*JcՉE������+��*��lt��𮤽'��.4E(�0U�w�Ϫ�r�N&�J��:Pͺ���\y�ڀeQ�9P�:�9+�4��DS��xA���qQe�XwDQ�(��v��@�j����-��F	�r5�r��B�t�����7�~Kk�Vg����i%��6�Q�AF}v��pW?[_�>*S�B�V���Jm��Z�R*1�ӧ��kWTt�z����mT�AOM�b�=_����W�1nZ�m�I�"�u���ʉ�0�EP����F�&�|W���������K����ȇ?�����E�����<C��NH�S�S��+�f*�I���wdq�|����٧�������\��_Um��f2�u1Q��2S;|�� ,�P�U������C���:}N���,�o.���k�2쩘��\Ad�T0Є@��+��%y��T>��O�U4�_��_�׮�uհ*4����5��s�=��X8�26�PW���3�{��Y3
�6`�T�=����[a��,G�W�����/</���<���k�ߔ��gA�\���{��4V�1�}���%�(�cj��_�%��o]Qw��䃟��|��W���׿(��������{�*��ܴ`z����ۯ��|�� ~���}��s�\�����j��2���\\M�1-�CKS�W��/~�W�a5'?��SY?���_�W�$����ϫ��;=RDB��8e��ӝ��^ Ϫ�P}X���UW�ԍ*�F��X��]��;{k�*��״�0�pB�+�J�{���u��j~�}@e�H#35�hS���L��o�*��SSwE&j֭���������??~�A�/�,t�;Cʾ���!�F-�������U?�����rq<����:�3C%���cU�A�1%����E<��wO���JEҹ�r��Y���t|�!�|����չv��a/��./`�A�ρ>�X=cP l�3<��Bew[U�N�������sO������8�h��N���d�RI�6��ܮ|��H�(<�?)�9Rք�>Pm��T%U��(��!�ѩ����j6����Ͽ|QzX���D��2�Y@��,mf�qq����Te����i�$T���)���>�A��st��60��`Z�8
,
SQ���.(���޼�;[����?tS�;��pX3��P��yaV'������to|O�d����ړ��A[���!���Q����2�᧰�Z+�,V3��4ׁ�j���-��J"=���q]�
Q���,�L�NTfF���HE��[˷��	�� b����������RY�h��4Q��pt����G�=������M+p��Tdo�b	ܓC-��K�0G��[��7��F���h�O'N�11יLm�1�?Pn/ʍ�EY(3"� �3���u�4ÁjX7j)J�f]szO.�n��ĭʆv�Jm䑊���w���Hmp�X*���t��*&�&��J�����J�!LI5;�rl�F�y$KXQʭ�+��*W�9��~�Muؒ��C8c�{b"V4_�hOVj��BLw�r||��椇��ZU�xA� B�O0�PF�>S�5R_�`6�RO*F^u �CZZC��}��DV��
�xkD��f��p|]�/�n�Z*Gb+�r�wƶma�����}�p����eO9&D�~[]�6UA 3�.���������1�ա����J(5\A�M�C$3���i�bL^��YJ����	6>4&P/��j����@��Q^W.��^�����(|�Ce��LT��؈�¯����1��0'�)��{�!�|u����a���%�߼'D**�u[�x�I����|��VBN��c�{`�C������jw���������=y1��ĲM�)���	�|��	��l9Iйӝ�F�@1��E[�����l���1�r1�|M	�.p����I�%�&.[��U1"�?���ˏF.��[l�9g�'΄^�b��7�
}����(��lċ�=�'���aĒ��H��_����8:=:���n�pt#=�<vX�a�a-G�Lt������I(Υ�3��J�JE�q�ql?\k��@�8��Tz����-i�υ������g!/]'��V���<�ם��=>0�![�F˯�����s�����)����)X��)�.�a6��+q��m� /��HXp=�
���Y	]�e�뙉�$�hk�8�¸���?&G����K~F��o��+R��}����Cp��6��r�&c;f����8����+�t�ӊ��pr�Ȝ%[p�׃�Ֆ
*QɈM�7���8>8P"��gY�����[��I��Y�|/���u!�����2���%��]�+�o3P^�m��³@Y�A1��ǒ�oІ{�ޱ����y�@h����v�?��n�HN���|� �k�q=IA`D�����i����	F�J��D%�cj��!�᷉�m�������|��V��r�Fr�O0�]��P�J}3�(wzv��r�o�`��� o3�$s���B����n1�1,��>���K[�ol�q�+�~,)/~^H�s:��d���M�'�����n�Cp�U�+���5�讒��D͘��Eo�����R!���FS�\w5�l�"hr��XyYr`�%@/�Vn˂�x��I��i-�Ct��%�A��0�f(��߁lX���$KpZ���f�`]�mȔU���#��X���A:��	�!!#$$p<T��"��&2a
�eh��}�HsR;���������`�T&����kP �L���F�$�8��Z��@*�����Gȅ`�֬,VpI*�B"AAޢ�4�N'd�
#8�ǎY���؜N]p`{R�L��`���dpzU�
�%D�bg���&-I=0�4ͪf�Ɔ��S}���n8̡�5�C��XKw�yw��w
���@#��$��}bf��>@x/�ˣ�.�ʵu�Ơ�A�ԑ��H�G��H�u�F�����ಋ�aa�V;��pgB�b~Gj ���2UI�5���U����lmQ)���e=�ٸ�|�L��{�}tW-e�􉮓0����,��+t(n�0G�n�6B�C9���h9E�HE�ޞ�Z��? ��mx��ֵ4��tJ�`9	bA�s:��(AR���{*��,ή��B�>���h1^|�
'|���&���K��f�b�d�r��y�w��QQ��].�2ra�� vyrsRܠ�x8������{�/�C]w;P�&"/�� �5@J:�aD��=��k�~�R��@��6����1֨��6�k~�QP"������a����P�~�$B��	��{Ő�D�+0i�W�9ww����������< (@SN�NNHx���m;3: 3�� �3
�u�δ�!�d%n�76����Ǡ@1q��J���vP���P6#klb����sr,�ХG��#��&��T����>,8�������Sk�1Q�vq5�oc��L�� H&�{��+���֚���<�U��f�uƐ���<K�~�����]�AC�[6��Ҫ� \�F���9F+&đV��|�0nb� ��6������''s�Z(Hd�c�Qۘ{���mK%U�g������.��L�@K�i"���ν|wpOJ�U�J�"$�s{Y�ъ{���lz�0#;��`,>�-NFD��h�4��ᖉX/kd����ԢN��u��zv���[���aV,��#,\YXD4���Z�oN�c�!J
�z�@�)��G邇Q �m�}���ݮ������e)&P`� &qf��@>��th�3U���.����0�-�+��
8XjS�3Ue�c��܎�M�䀦"Kd��M w��.A~�,��Z��0W���"a ��l�} o��F��>~�9bu�I�)D-��z�M:壻S��v|�(�U���jz��v(����\zp�"#Y�i� r�1G ��z�h:�%Qj	�9�F'G��r#a�*��#>ʰL��Ȭ*|nH�S/(C`A �;c&��h�(Ԗ^s5�s,>ŋ"	<��Ň(S�=Nc�T����Ȍ�������J�0�t}�ƥd|zO���� N���@.B15H��U8��b䌒3�Q��J��2�������ۥ�3���@��ݤ���YA�r	��r'���R2Hr� JӁ��4Qg��M&;�0��#z_5��pj�O�6&΢QMԝz!ce�f\�I,��a�ߓ�Õ�,�AY��	��
+�B4�R���H3���jCƋ��_���0��#��3yM�4 b�P<��� $`�a�к��\U��˝GS��qx��p�9a�f,tfU�<7��d)�?;�M�;��!uU�����b�Q���+���D��hK���
��\�v�q�6VY�8K!}^��a�1H�t��@���= RHn'7�ĈGv�IV(����W�޶#�|Ki�bI���$���]w/�����tb5�4bL�ʔ?�.��d�}�1P�\�t4��b�V�C�kVy�����c�����N��� �OK�3r�Õ���@0[�Y��V���D-Jle�˝���@������V�QzS/x���f9�<�eum�䖏�c��0��h��\���5W��*�Dn7QX
��~��q۸0�)'?�_��&�Z�bO���3k���>��-�`g���'��;�g �Z��Z��ڭE�,�DA�n��֢E(�/V&��<�����cg�S��Xpш�9ä�!���xa�)���d�"���X�l$��Q$VV��@����r���`�E�"L���%�Vډa�	u�ͬg�n��G���Li��0�|1iJ�Ո\8�'���a#.�}/�m:j|v�kT�bwn��O�0qb�>.4�ض��\oKx˹�H��A�S|s,)`�k��h�)�j"��<,�of*;WK17��β@!�����̾���T�b�hfz���;�	0Ya���Z��
u��ˣB�1?<b\>����Ib+j"7�,3baE�T�v�=1R:�m1�Ep9VU���t/��	�LLo�y�',:;y�9�c2X�9P�����踕�ru}8��x��R�%�`�@�N*YO&��b�� ���`+s�bpXX����4���=H�z���fT��w�=�ݝZ�۠t6fȖX�z���ܛ�L7ݤv]�x�y�oZO�0q[\?��9/���sJ��1��S�R���>c�-z��.<\���	�����хAu��w0���QQMXgKj�����9�l�PT�����#���]R�wZ'�a�+��ޞ
���&�i�x2��Gɖh{�%{�w�1NJ�G�D�24g��K�,
��I�v�g;Y��3;k[+���E����p_h���;a���#B��mhN��DZ�2u�J1ڹ��9l��R!l^����a�%ND�����Ќ�%�3ci���G�yXULV��h)���@����߄�%@��eTߋ}�.>�G=��	�G $��s!��\���:�
}��̑h���-�ROw�GpQ��-�� �N���	�k#���r���|s+Â|6AX37	��1���ڪ\����q�t�8=uȴ1�F��7�,��9 2yE	���u�т�Of1e���	�߄��8B�nE��z�56:t�{	�{�,2nmse3����]����Y���U�,��u,�@��i�F]R
�O>�9tט<�Шha�d��{�,�P8KW��O��}8{3�ۯ��n9�����d�'��Ž��cٚD�pP��zɢ�JM?�΁�o.�f����H/4�F'x�Z&�W�B�Du�v?�`RZV���ؐ�e��	�t�� <�͸,�����!��M��s�6,�\S
w�8�"��`�dA�K� Y�>"��� ��x<V�ʌXȖv~;�g�,�V�¡�>����,�9R«�@��*	��&��#���.Nu�)Z4��c��BÍ8�X���3+s�6�On��$������F�/9�yC�v`f$e/q���}[�=B����d���,�?A�R�{Ö^���B��$T�/k�^���IT�DU���F�������� '̖(��6��U��$��Lv�Gg�d#r
���v�{ZC'�G�y��2�o��B��	�&�T]'�5��$.��9r2p�C����˦6i2�?�vx����^����(e�{�#����s�y�q�����d�㒈��:�B�1� �fᒋ(�2l�"�cM�g]k���:��,Jx2�wM��E�0s����e���0�Ye�|��[��|r�cI��SU�L��pe��׻�0��3��#׋��G������:�[�n��y��Q_�b5b�����*��*���	��}w�8���p؊��k��������V��lp�}��߲�gqGl�<^ߵن�b����H_^�<�$�S(}���q���2qlN����[,��8��]]��N�L(zH�Υ�S[?2;�T�~,��{��I���3���>Xq˛�(c��?m��e�X��D[VKj��󯡪n���9�u�%N���Ot�4�-Vp.1l�E��R��Dw���N۰� �egM����2��9�1�K�)�P^����m\�����zº"��S��Unc�蘐e�\Iՙ�]�Y���;E��a�-�N�($�7B��d�'Q ���q�K�	��Z��х~e?3�g� %ژc��7ߞ��&��b��F��:Z�\;��St0��~��V���X�ƌ.�ҙ"k���-K��M6�?�P�Q��l�e.��B�L\��új���oD"Ϡ���s���JF�u.�++%�9� ��h���U#���G�e��W 8d�~kz����x/�ɢ2�?������C�(�T,�����[v��P���to�X����T.�o�/�[n\��A����P�41�A$A�|)�C�ܯ��tA���=p�Id�V@�-��0E_�#��+^邟�ϝ9�JX���J&�1��9s�-x�a�J72S�/G2B�����+�NJx3�"�4t�Qj`��oK�m���斣�o�ܚi7���t 4»�>o@�9����/����/3n�	+���@=\X�p�@�<�f�MK�~� ����I#�O��A��M`1�j�0t6��	E#����8A?5�yM�����d�;�a�b���&S�۱��
�f��ypa��.�N0/Ъ�+�%� d�]$8�	t��5�)B��+Ƚ >�1�Uwf�8h���eaT2	�z�)x	�xE���h-S7F4̩T���j�ɴe$���;��*��	�u}cowj*�5l�����l���s�N�OG��2����#���ј2�y���ã�X�C�`���l�N�x,	Vjd	�����{]�a�k�2 �t՘��x|�{@!� X`T4��r l��'
�����sb ( n���0A���w��p벐���<���xT���oJ>-9p����y)���7�a� ׶�iWt[z;��mWS��kF�w��\8�,��,׋߁�R:�$j��t��`������E
�p���<��LB*X�?_�׽Q#�[h�PV;��%��� F̞48�ʳ�Vk�X�~=bh���G���J��Aa�7�k_ a�O@Kh�G똔�М��Q��jv��2 ��x"����ղ����ǞU��2;� ���Q��w��NfN�l�8G�a��Įy���}ۄ��[ V�X�}e4���D�h@���N�0*��7q{�͔�Xk�h��H�\�4���Z�3�;B܅J���:p�Q�B	H���{��rr^ȵ���r'�s�A��6�����R��QOߣa��j���W�6�m^4�A��tÒ����Vb�tf��w%��T)�����A*f��)�]��<U+s����Q�J����01�'�У7�;@i���a�v�2i�3��g�M.�^*�$�h�������Ȩ�����Fmv��a��2<l��6ұxGЎ����e�tK�iYR�.���#�=Ũb��]=aˎG���J
�!�u'D]B)�!|���h�X6��7.����(]���ø"���%��2�����*�Q��EƎ��o�Ü�����(@��(F���3hT�0AW��U�T��_Y��^���z'(�l�؀�^;`
jI=����w�qg;��7��"Y�b�r���2��Q��h�?ϸ�k�a#����w��*=b9l��"pl����e��B�u�41��s��.��Y��B���$-*1��G7���@�e%��_��+TSd ����$ngӀh0��R._q����0��$�R�@Q[�.mp�x�!C��1.��=TK��dk��+�P�ˀvш+l�
�ebg��-<�m�$@�W)3�l�8g���.B�96A~O8[�,�����gl��K��}r�߳�Xr2*X�C��5��8rk�Y��x}U�d=g�`=,��esN��-6��J	�n�W�M�v��}�4���ܓ��t�3��]�0�"���nG�B�ַTY�q��V��a�@��`�1$���~@������B`�x�G�l3.0��,�B2T�{�.S�1�M���%X�K<�jܖ�J���XE_`M��	�d�k�Sbv��.��
���neU�F�������.ae:LpG8���˃i���C?x:9��gX0C��3��6���"����?҇-`���~W��%��b���E(F��h�EgX�jU��#͊�N�V���e�b��B����W׭ܶ}���)��a��������ż���J���>s��Wli��?0���xn�`�o�{�����eJ�\C8:u-9��L�2a��
�|�x��L��l&���Kff衑�!���Rr��[/Y\?r��bf�]��@�y�h�GR.�,ʤh���v|�ǒSAd��I���w��+Ļ=�"�g� �J;+�a��5��7UL��dc}	��Lc%|Yr�wA�r�Σ��,-��GM�Y��:����o�رi���8u�[�����G<3"��g����d���zf��O��څ�`�7�__E�S<1�Jy�Mܚ����h�>8��c-�gE�fc�����r�|�b�k�v(����q8B��ĺ&�q��\�6I��	���H��T��z�rNQ���vY���E�R�g��=3Wά�AD����.AɎ��X�%�����B4�PƓ���1�\��9�c�3���(���*��NB�X��.��(�@� �Z��!x9��t�b��l�f��he��� �P���g��f/r1Q�y���òb�X��B��q;z�[���X-Ӆ�,ܬ��,R�Ʋ"�KUǄ
�w (�r̒�����yX�����2�0�V6�u�{`��	>��~�d��Ea�vqt3��ɂ��xl9,�(�� �"�$���i��	���F��Z�5U�@��0K�9)�$��޸��΀���J�Ύ����ɲS"�̦r���Q�x0-��R5-����`�K^�q��j��	(�i�f2~�_惶ȑ�B��oJO>�ɄfvP+����.ͪI��$��錴�Гm���䛊��[��[��"��ڭ�.|�Yx�u^n)��(�*��+#
ۥm�hl���w�!&�����ʇ����x�w��|1&	�]��Nt4�D{�����~�0 '�J?Y��*.g��K�U��̲6�!�0�dA�a��v�"�!"~�}_1����)���y���L�DY;
���_ܺS�br߾*9+�Cp��۩�^G�B:x��ob$N�P�I��X��� �O�-��e�yr ���i&2�<8��`wjI��<L���@��!=�\�)^����Έ��r���8��j9��?93�*U��X�&��&G��B7x�T��ĭ / f�#�ES˪��+�î ˁ�>��v��d�����;T���Cȿ��0yv\����2����� {N�Q,���HA�
��
��\��^an�0Le�ˊ�g*E��E�	�(�����H-�b��h����ӣ�>*贱`�mخ�B�|�X�cDe�f8D`)FhF�-`e+5Kw8c'���h��pG�`H��S����/��ְ�=���%|�|�y�M�̰�dDg����o|,V��
>�4nP.����X��e��2��z��6��_��k�-O�o�(�qӊeU/���w�bz�s���lW,͵��]����=rc	�
�nB����������$��;���60�"��%�� 2MG�4SO�Tq0�wV�<�vM��Ɋdr��		����bZ&
�n�		���o�ڭ�V�$��r[;r�M�Y�h��K�yWc"-�+2��v��	cEx���q �İ���yMq¤]�Az�������(.j���R�o:�Ln5�*(���jt؁�i�����U��A��ћ�� ���Y�#���q<"��|-�S�+�ܶDz����]�E��W����)�ά#m���C����"Ӗ\��m��4�OӮΒ����-Z���]�e�܋��qp��o �pM̥��#x�IB�C��P��C�*�r�"94�f�El���6�79v�҅�Ky��75VV�g��Z:���׭��&���&����!���ˎ��Y�>�wrQ��,�����Q���b�l��I���(x���Ak�H�Eg�]X���4B2%IdV���IF
94��}-LLGb��� RR����H�`� �f���2Q���%�W�;���^Tm_ᤝV2Ȯ�v�[�V)Z�~m�8��\�����JnT\��	<�<W���Y��V9�l�:bH�w�����5|(��_�_'k��\�}:�xG�&N��13��
y��d�q���bȐq1�;���2�]a<��}�K������z�ԣ�,θ
�Y�|6���Le���k�_�ŉ*��X&�.�Νs8��A���be��:�VB�j(թ]ZY9���R�����d�3��EP��DF��g�l��Q��bzӷ�����_�M'5ԝ��ER%�
��:�=�۾4_E��a��H��x%r�XU�z�k=4 ���ݎ������!�L?�X�J���:��匭[�.�_�V�@�hu����8-�ޔju�C�X��]���.���-V�iQ��-�8�����~�٘3O&�L�n� w�[o�
� �m�cJq,�L�~b��h:�\]��<>�*2��x�ag�.�ǉ9����ú��y���h�N�wґ�d�΂�ڰ�I9���d~q�4�[f}�m�6n����$�U�ա�q[[�'��}#ά�V�ӹ-_��>@+-j�nإ5��齃�4�`�P�u�J�0#<��Y%�Z�	2�)jk�a�1?�����L�Gh�_q�U�9<�"��Б\�M1ԅ�.�Z͡`OCg_$z�5�����@xP�2�B�vjo��̿XD��+9�*���ῖ��sB,��-q��7�����Dy�Ie�'FMF7m6=t����*��`�M�
*��a_6����]ʖ�[udn��-I���Mr9#��daηH�܉.����+�J;��9ږXȐ�U�IwJ\^gEE�fc�4���(�?�(X�ѭ��!���ʹ4��E��l�ׁ������&r��w�3���^�lF�f���zG�jrN�-o &��ګ �ǌ��ݐ�(������~V�����Zw���\enD����C��Dx;r4�<T��B�N�@��WW�DìJ�D)빶�S���C����d@�鵷��}*N�e���\d��Y��6�Xv�;e�����P�����bc`UJo",RhU����xW�dB���J�q�8g��q��^2�]�\��ԔeA����E';��-&�6hJi�3���m��pO3]䭂���)�tө�]��~P>�i��]F�
9s�;U�Fd:N�.
��|D.�T�F(�1������\�4<S�=Q+T�ȣj`U$��&�呼(6U��"��"1l��[sN����KXx��>oy�[�l"����-E�l[x�RSZ�\�kv-ȩ[u�=��t���>�Bd����u�L5L��yR�`H�fDv����l,-\�\�4�q��a.p|&�47�C�	ɻ��{9�2��N�W,ۍv�Z$�Ds *{wV),e_�+��mѲ1��膇8w�y��9!v^ag�AP�ۉ�2X�1'�3�3k���p�`ֶ��D�#N�Fq�0�D5���1h{�s�E��V!�C�ܻ��(������.�S�բ19k��� C�e�{�k8?�"Db�л63��c��n�Z�[�[ݵ���݈�-�j�)"�ٺIF�D�{����B��N����L軉�;utz���'���m�Y��������Q8q$#�����""ٮ�n���qR�$�T��C�&��[GL 7k�����m�	��Dr,�,���_[��ޔkz_`��ם.j�dS՟<�f�PdPj���D�N
)�7-lЙ�ø�B���L�h+[�`�>,��i��i1�h(c�.�~��b���|��9y/9�M���~O<�3���M���5��=x)Z"�Ȱʎ�K5=����|)~ �'ѭCj����M���U��΂��+[)��P����O��A�e��vS�s����R��{����8��L#����cX��̢�٤�*@p��z�� ��z���ɘv�2ؙ�`X�9W;�H�?���֩	mY1�>���St�2�';�č��N;W�L�7Ȇ0��g�}
o��6�;y��^����Gy���޾�<]���=���D����<V�P�	(Y�w��tx�+��l�����#�<p%��dmDuJ�dʍ��N[�ŤI �mv�����9� �^���nN(j�|G܎+��nx��V�������#*WI&eɾH����(�Df�������k�� �BD}����W�ƅr��hz��Hm��~J��-V��=���W�[�8.�#*���ᄢ�h�R����%��7��V�$��[�b�v�5��~�oY�\Xv �&��]�S[?�L��B�)�hE0l{���@��ꯨ c��'����w��7,�/X��qW�JL�V�8���ؖ}��W>���t����s]�b����v�s�k�p܉�n;�s$ B���Z$�P��<�["0h���>f�cE���yپ\2���&�i@� ���O������_�#���]α�ޒ�<�ΠC�����ݔC����T(��j#{c��?1�u��P2�&9Y�ؙ��R��4{��<�е�_��.�Lkck�mU�T�7G�|Kş���r�=�����'�@����%��z�����q1�cJ�O}�����[td��#�V�vc,�ɔ�Ȉ�!��>�Bb���@������A�q�X��f�`2r��jp<� ��1��2H���m��"T̘�iß��]�����9��������\��%��l�dIͤ������5>��p�{�1����u�G�5��#�O@x\ʥ)opu��<���N4@��x�0� ����L�k�]�N'�53��v��	ָ�s�0w�+�.�� �̀�f`<?t��6/�M�G
|�lz2I��dX�,7��[�^`��`.�6�����!vw������m���,h�ab:9�#���9��2�<��är�/��VV�C�x��M�C���"@�d�%�s�*�^��u�H0��։�>�<E���Ax��=lZ�9lNOF����D6/�H�I����rҽ+6����C���wo,�Σ@�4�ͦ\}˨0����"9� Z����/�L�E���� ����cW�����Kn��cn�Z�"�ɚC$�A�w���f�l"̮!��tژ�v[��؅k�K�o��d�O@��F�Iz佢�d����(X�\[�Ε�&k��Y��"J섙�h�N��Z��z%�6�lW��+�M,��"��VN^S�[�%8�4	�;�'� �	�M��Mض1v,�n�WEmG�a��*��3my��P�:Ή2��U+5
����.u��&��k�IU72R�q�D�c%�PKa��P'қ]�V]�:1��1@�,�5
��āo���ȇ���"�{�O��Xe�p�@0��;�@�����߭�G|���Q���]�Z�n8.�LM-�uc�0��m�����=��Ӓ����*c���:�k�|���wCx��b��JdW�����K}�a�wp}�g&��b����f���v�d�S�iBOI8O(T����b���r��	�!ܣ��@��|!˃ci�IZH8S
%2�	��\�|U�ျ xIx�ƥŚ�k:�.�Uu �~]��B���oV� ��Ѝ[;���mk��z5�^����#�p�0k�Q��w<���U�o(��!B�#��-����\�6\��`
����v��ߏ�P���?n�[u�c5@':Ik�'%�2Z;A��2���}�@)G[0�1�ɓ���֚1ԅ�8�����mW/AԬ]t��7���й',vD�I	O[8�J%�Գ<����
�Yu�x�:��+R1���+��P*9.�N&"�p���j��֠`uwY���`]�fi�14�ѿ���0�Td�7�`��v�S��*��c��/s�^b+�7|���V��'#k����$Z7�}Ψ��Jʢ,O��8_�k��e%LQ�2\�d�T�⨄�3�=�ſ!|�r?/+3�P���%��i��$b�e��u˖�ּ�
���>1zn�[S[g�ά�ܦ��㜷S� h��*�:ݦЁ$uο5��}�aP��(c�x1�G��Ѣ�^�ݣA���k؉��J��s6�vt��z������'���]����'��{抖�N�5����+k���T��4��q�hL�ZVX7�)J﹙�&�2���d��]f\���-��y���-;5!>����C2N��Iҭ�Z.b��8�4׬4,Q�Ү/rۨ����	�����6�yz��g��ڼް��fHs�.Ő|��m'#��89G'9�#v�^�*���p��Z���/s74�f�����HӰцl�`�Q2�%�`{As�� �yEۚCU��]O}����aQu1ډ��m蠰�ۄ�v�Vn⟓ȹ�����a�"l�}ͥ�&g;����Քm���<|�}r��9펙"Dt�hv,�o�՛7�����[z��v��M?���ț:�'g�v�U��"���i��E�e�,z�Ƣ!���R�j��LƷֳ�m�B�Xl-QZ@2��E�qY�([@���2��l��3)�M5o����F}xM����<,��A9�� X�m����SCy��GeV?(��y]^���\�r]�����Έ㔫���D,6��z�S�6Z=y�&Y=z�ĺ���!���u�:�Vg��(XL��έƙI��J��1b�Pz,"VSTlY�^+��JR섁C�AF*��򖧔� �z%�NMe~��7)�G?��<��i��rj���/�{ge��.���z�M�`f���rz�>yq2��rI����Fw��d���ʐ\�XO#븃M�~�Z����#�j[�Ě���j+�v�Ӛ۹N���w�W�:.Y�)o���?���L��L���Q��Z�q(+ג��7ԙYUC�Ը����Se|I1c��u�,o�ٽ�|����Y%����#���O|���O�):1�V�z]�ׯ]�/��o�|���}�	B���M58������]
/؎�NV"�r}���K4L5k�5�}���iK<����[��N���wO��+�)��4n�T*G��ӋC�ouS�.˙�\�uT�0d���)Q/����S���iY�㕟�I�D������&���o����K}�������g���?*���G����~|�u+QF*J8�'���N�7��=y��<���Py�ڥ�$�!7Jڲm��L߄�څ8����J���Y�+���P�ϓ��~�Hn��n	ߖ�-^Z�JR�e�_��b��uy�芼vY�-dG��1vC�n�N�P��f���\��oĉ�G�ЦϠ��;7Y�����+����������H>����՚D��Tj�a���,���O�^�w_�G<'��s�q�,����V��0v�n�j�Λ!��#���1�!�����cluS�ʗ�	�d�Bn_�5jrN��k��壋krvyC�Z�]J�y�ّ�Nx*#U����b�zu���X
��eeg��VT���=*���2-�*^>,ݷV�
��%U��\��MX���ާ"陧������Z@oޜ[���xD�\����|�I�=Ҏ~��Ys��rt�������'�Cl�ؾ����}�^���7�jq<�D�[X��d	�����K��Rf�T^����T������t�y, ��=��}�U�.����Sc�r���*�[tOBC7q#�kU�ν���#O?./�YNM�rn���r{�f>+�K�{�V��I;E��CF����?'���lG{���*����5� �����Œ]���#��]�3*VS�>�2v�5��������%vd-�y`q,��CUƧ�X-����;��� �*���Hv'8�b&�S��*p�����9Ƣ0���%��П�1L�=�7��ّ쫒f\>���c;`֓��
�x�e��NM�����C�wT��2�������;�}Y���v��8"����iyw����6����r议�)%j�����;�l��4�V-%�d廢��`��8����������x�PM��@k=��Xlo#���D}6�` �'!ptw����Ǧ�b���Z���8~Ӆ9���{dq|U���oȥ�Z`����⫯�O�b��`Q��:��S2��^�O�����N�gHy������[�N��'�l�*�7��R��e%6�G����L�S24N�1��%�gJ�n8�q���|�8$``�>�.����J��X�N��y�=����AW��Wa@���H�����d��̡*顬�)�������6:�[�}�{����pd�>��/N�9�
rU��Y��f���81H_V��
Y��x#	�V�ن`N,C;ZX��Rf���&%��� (�bd�p0nUz��+��C�7?���vy0�\}��.�N/cG����5�2�2��dﴷ;:����ysH�NS���b�v\}k�^׽EMWX����d@��j�6���fT=á�X�is�2䨜������tS/���E�X��2��Y�99o>_���L<u���ƛ�~�T��pX�PQ��F�-*�8OH��/�.G�H)��54�F���7���X�V�t���\��z�5t��Z�^���g2Њ�ڪ a8��d���2�l�3W�휖�r.St�f��*:-I�Sn��k�=ym�/���ZsnM�>1�M	�#�~�?REэ��N�A���5��?���6�R��(J���q:���r!ce��/�*�u'��s�h��^�
::���9L��L�goWy@ T��ǽ�m��nh���h{�~5E��%��תPU�\P��7��!Z �v�!�+�LTV��9#�<}�|g�\��ʑ�Ȇ@(L�rH���-����ɣ��Wo��7oȃ��<����xP���]������?��f�Z4������Z.^�(��ղ�g���֍\֍��;+�MǨ�ݥ�8k
��
5�\�tc���n�����Nš�.,�V��AH M�L$r�;�:��=Q���oT#��J�s���)]�	��(��w�b��$p��cZ�s\�~(/�t^����K�廣R�����%������m�9=/�����o����I.]���.�����T���t
�ϯ)��MG�ޛeC$`lbAi��c�:�� �-�+s�n���Ȱ�qΨ")Q3S�YM��u$Gꬼ�3U�(b;Ki��!����X�O�䪊�U�mGa1x�Uy@j�o�)LG@i^��&�~v'���,G�����~�1�ݝ=��E��k����;/��9Xv2�]�^���rniݵ����x��4�<i�&�*��8�8+u�%��<ua%��fz�ž�
�{;P1ƕe�<�E_�+/�Կ/�&�� �  D�B]�y��e9f��N���>��ف(��(�>C��?[ȿ��s�~@Ə=(�/\����<���d��C��@Օ+��P���B�5@�;��$����V��[--�2,�>���Jn�b�DfC0J�C��̨�R�d'K�C�v�����u��m�{N��ݣ���9�m�q6�t�hU�.C�
���6��l��&�ɭ��F>��Y�$��hĸ�JM=�h���`��J��Ǌ�H���[�W����v�M���ԺQ���7����X�=�f_�v��o�7���\[�rШ�G<�r�ƣJ<�:��/#�8����{��F�R�"��<�BU����_F�m�y1���T^>n�X�&�_x������V�iǧ�j����Y���z������<&�1J�a�^�CU�+:(���8�&#����F����X�vF�廯_�7�U�|�!9{z_
Uԃ�>O��|�������p�K�*��ឬQƃ���Co���J��S�TMb����؞1BI��Y-���g��_��N�W���,嗾�=��ﾩ��`�!qK����?'"�lv�[5��z�F��h��1�H��̎����豣�{�*�C}��`���a0a�a�S����= ��T.]y]n��}�f|�P �X��옋>�찂���lƄ8�I��Jul�.����f�~�U�kS��u7�/W��8ݸ�r�����L��vsJo��Ԍ1��ポ/�����<G�xH-^��1+��L	2��i*�D��r�V'i.��7݌rjoW�a}?�� xD���ҕ��9��a�~r���j)�T���p�Kd�TwJ���c�������!��C�.,��Cuh��VH�����g��]��l�T.\]�'0��6_�~�܎������e[,Cj���h|�'x���U�ݔ�r>w��*�������am�F�o�H�nD��)����9�*���g�vwd�{�fb�C��4�C��x6j� c�X?�o�Og��3���kQ�X�7<B�]=t\�{j\��k�б-h�/P���&�Y+���v�����>�V�����A����ngDmnq��U�|�6;>��s;j"Ѫ����b���o^��w�)�1Ӏ�[bw-uJ��O0W.�b�*� N����[(�jdV��rA���Z�g"�^����P����6;<�"b��Vɩ}���7�d kJv�)ke���K˻���g������d�Er�F���;����*H����'�/��3z]�zM�I-�z!g��(QU"���\^Pw0ڧ�;�ӟ��^�g\�W_}U�J��\�xQ>�̳�lw������b��ޔ��	-��Z3z����|���SO������O�c�=)_��eg��<��g��͛긽��8������J�ğ��2)��^�v�ʯ?�����Iӱ#�t���&e�
�������H��u=a�~'��[4/�v"A,_��]ʃJ����>U�y�7C>�#��G�Y��� �{�C��#�2�}������۸��׮�3zV����r|�M9T����?����l)���y��}�S�?���^�]</�/�y9\6���������xn�n�g?�	Yݔ�j���?�G�_���ď����~E�z�9��g~T��{�o~�KLr��//�b*�?�Q95�+'��KWԑj� n�6[��srw���s��>��j��(��?h�jF���,�y�{�u�v��{\�~���������E����d��\z��s?�s�S?��(w>(_��2D�����#���_��_���?�Ay��o��OX�i!���/�g?��ҿ�'������ܼ~ ��c���-)�.���|�O�·��7_;/�x�i��/��|��?��)��_�翡V+��N[w�V�Ҳ����)�ME���g����jZ�'��w����T�"'��n7mF�A�����2���v�����0��?����^�o���?�q����������a�.r)��P�|�j���'����z�If�Ν}���=��g�ܙ��s��>&�����P���r^~�gT~쓟��������ß��3�e2��5��x��I��V���TQ��p�������W�o
e���d0}\��85�����g�H�w�D���hP_�#ۥ��%Qe9=+��Uy⩏ȏ��?,/�q(׎����������gd�s�|�sP޼rC._=Ro���t_F�}����\�vhU�E����?(K�&�y妄��������7y����99u�=d��_�pA~���r����?xEv�{^���q�/ϝ��z���*�������_��|���`؎*�v����I���LtA�z�;�h�2�П?{'��߾��y�������0k0P��"�
8j��I\?Z�?���(�������/��5�e?��UV��Pa�r��y���s�H��E��?��n�yY��9C �x���ټ�����+��+�گ?/o\z�%��h;:���ã#�@F��/��|�׾Ά_�җ����̤����<��K򘊯�7��S�t�qT6��;���[��,Vs���Iԋ��=��a_������voߵoc�ZR؈_z1��GX�=f�do�'7���j���/��{CUd��1O���=x�Z�Ǉj{��U���!F?���r��i1Qb_������^M�W_��Ě��cO���7���N��>���U����gO��b&���9�߁^eC�M��_72@x��
g�[�.�>[�dto�\��_K��?���W�wp� .��e|!��G�7�̓�r�Ԯ^�&ו����3'2�%7G*3�*��c%zO��UVr�VMZϙo�B_�U5�ܶ��tF>oOEL�'�,��xCMĠϙ�G�ڵ7I��gU�TT���HE�Z5��ǲV��O�P��G�mq�PcA���O1��|�*f�����wJ�{<���*ض��Z��������J��߼fEe�]�*z���zv������g��}Rv꺫�������K�����ng�f��ae܌�~J9zS��G��x�~���K��\����fR�*-uw]|)Rl�y8����ꎰ������[p�z��]ݹ�H�d}��1�w��n�|q[���v�A�#KC.eIv��j�]~�Y]zE�P��0.j,�X�,ܪ�7�����\]�b_e)��^!��]��q��S�E�G(Z+b�5�4'�En�.7uw�Ï��u�v,���<�pe�ߧҴ�"�2��avK�x~-�����{�E�z���֪�n����C�ecxz���S5wB�*?���0HF��r&J���G�' 	��^�kUn���"Wt�TNV�L-n(Ӣ�]m$���CI$;g��B��b���'O<¿\S�qz��y�!ځ^����������<�E���4!O��� ��r���Ee{���j(+]�+�Ʋ����U����x9�ѯ�K��@g@�s���=/ŉ�d�VÕmW�:,I��ܲ$ٷ�)�����r[Z��T¦�x�_��k_%�>�Z����[�(�z�$~��C����ÿʒ(��{�ɍF�Hb�M��� ����<���9�5�-�N������}Nv����/]]�k���y�J����=�����@d�r���N:*D�;A䂸ET�K�U T� f�	m�x�|���gA5vb��G|E/�Y��U�����3�ʍr�8�<����\�|��k�㤮
~���Ɓ~'fI���F+C<}�_�{�����@��v��^��wF����l�ڑ�0+�?�dEd���<� �+��PZ[Y��Dhk���+��Kd!�Nԏ6�qu���l ����S�ډ��1M���Ί�ge ��H96���	%�ϰ��
 >���޵��u^��g�˜��s�=��61)6$M��Z���R�����_��4o$��<P�$����}#B�T4��N�_�:���ˌ�s9�}��g}k��̸�N�����h2�������k�o}k8�Ҁ��:F}`|~�(���VF��@QĹ_>{ݽl.��u���ok��]�w���"R�!��H�r#��R$t�n9�
]X�d��Q>BO��{�]��-%�%��(F*��M@x
A7It��-�h��)D�}������/�ǩ*��M5 ߗ��5�.�>\8_���/c2�al���P; -5��)A���9]��	�L(������Ǐ����|�́��[\;����џ�QD�=�횙�\���*�}�{�*@���R䚕3o��:IT�מ�85�l��S/эפ��!i��u�.w*t��7��R7�1Brk|���sV$+[��&wv���>�®��ߥ�e\;��}B���Aj+�(�U(�`j}A��JZ�o�#����O������u��R,�'�K�Bg�xzpB7+d�՚���~���/R��<�˗���cCT���H%�V��a,>1E���H��۷nѵ7����TU�G %	��.j~}�Vi�����>??�0�7GSt�����,�½W��Rq�=�M�,�w�V�%����R�T�K�"�+9�kl�~��*Ҡ'F���-���7]e# (j�۴��,��.�x+�[햦V����T����쫻5߼y�q� 7���T�U��af*P�C�Pg��L�	�U!�Vw<���%���yỻ�Ԉ�Y)�[�1D���t������ v�>�w1�.+Ͼ���J�+ש�mѠӖ��LK֮��xH����\�Em�N��o���+�3jq��J�'�(T�.|v�&M��A�^�N��cs��s ����,q���9�K��s��d�3% K5?e�e�&+89\��T�اj��D`FW����t�=�(!�$�K˹����!�l�D�u��	�H��qnu��Y��msT�7)�����8��'��A���s�����6���lҁ�io�:k|P�Z����n*P���P�\�0#m{eP8�z���Vg�Sf��o���Ǘ�eF?U^*��FG���"pT� �a.�/v+�5'〔ȉoq`wG4k�2mkM�C=�\����[�5~��?f�T�@�0��&���1�*�%c�٠N!o�5h����}���:�_�B�ܗ��[l�h��u�zT�kF��ݻ�q{P�B,��cI�/Ǳ�o�U���{��-^�E4�� �^P�ݔ�R�f1�°$T�XvEA��O����9����k���a!�%�j����HL�}P\�I+g��x}�4cop���ϡ�w3��п�(T�eڢOAL~cZ �hh�1�eǕ%P�W�.���ƞ���3�jx�g[��ԝ�2Y�]Y��bz��Of�>��T�6n\%�s��6�_z�s��|�	^YQ$�EΪ1����!�_�B�|�nm�3�0��	�����
�4�h�����t��+����� ѢM�`w�I.h8A�ϝ@�R�2��4�,<D��=��õ�Er���+��)�
�E6�PM��ܸq�+�X����s6�9�R�mC�>��e7h@w�������Zk�Dv��2E���6l,��hc�!~���gM������)��;O8U
6n����t@���8�)�Trmz�/t����ۜ���=���8���`�Z��M�C52�en��>F���o���k�����hbn�!dC��
'�`���"DbP&��M���㖭@H29y>�T\]����V����04�Zc�g�i5�d6Ne"���^�ϴ(TL�T���q^�Ż?D�F���8Br����V]���{�RD�A�",���)g�������-�M��5��I����p�V��k����UF.~��@֩û�T&h|� �ɍ��L3C䚻�p26�j�璁E�-+E/\��<��=WS��Z�~W�9��e��v~�Do Wzv P�^L�.�С�d[]��th�üXy��Ð����y���i̻���@���u�j�И�:	U��N� �F��gL�t��:���QW��;2t��H�ʁO5��n�w[ +*AS�p]҂��F�6E�'FUeY$�ʩݎ�@� f2���a��������{�@1HE��/kD��{i��nRXm�`D?H%= F����V���U=�xbx_�12�nN�����} 7ؔ2_�ςJ\�z%f�9�C�f{�*���H8���t��`=�	An���,�Ui,�H!k0H� �TMvQ���0L�h�yg���E~���K�INɠ�
���U�v��<���ӃY\EQ�OS!�L38BZ��Kkk�)s{Wï��[WWWV���9���<AG����.�c�T��QKyyȠ�X��r��ic��w.\���C�y��0}���TM��8vԇ9G���Q�#U�����_��J~H��دҮ�9�e�Zv��aB1
�2c.E�{�t�<ml�Q�Y�G�?BSӻ�,�k�������
M�ʁD6'���Θ_ZO��ٛ��qG(��qW�W/���"��7�Jm�|�[_<4�[�{�pjf�q�'&4]��z��c�l�J��cJ�?�[:�]���+:����/���6!���6�e4�`߂ 1��z�<%k��	[�#Gf��������W)E�M)P2zB��%M�}�e~�kT�]���)ZX���I	���^�H�O?T��Y��C!��dH�=�ǂ��F?��o��p�fۻ�҉�7N����o�r�w?�Ks�)�l�����itc�;��]�.4jh�ms�G�_#�hQ#��(k�7Z0.}� E3�q�� ���U�jrH6܄�tJ����@���G"�D�g:V�W���`���%�Gv8� م��A�¹���PY��Jy�j��`�����������/�x��s_{��0<��N�h�>���]��=�{�7��O�N��� \b���"h�F�BG[�tW�~7�l�M-��	���؞U~B>�؈�7)<�Ɍ�S�2�y�u�*y�1F;�(�1毲��s�#%G�V��M��ª��|����V3�/�|8F���k����_���$YۯD���**o�4�������e�A�|:!qɭ^g�핕s�/_y��~�<}�?F鏯��}v��g��x���n<Y�F�^��O��H��+(��/��qs��9EȎ=�T�L���џ9�SO>�t���s�02b��$�%��݆Y"���:o�42��$Ju|Ȣ�I*��uDW�����Ũ�Wr|l�ErF=���*� ������[o|�ԩ����z�k^��c�y�y^����c8�/��"E�%�s���W���K'>�Ч?}W��S����l�����c��݅f�W>�},@ �g43�d8n^�3��	��P���J:ZT.����]��'_�}�YB㘌�e<ak�﵉j�Jasԁ{i��N�ǔϳ�@�w��n��;o�$/��g�B���	M?�՘��?�Q|B�D�eȇdH �U�lK
ַs���3U��:����N��̠�Ky�}C�,�LJ����6~�:��x(�/�~�KEPb�tU�^ͤ�1������/��}�jvW4 S���~舆n���T��瑞eк/��=������	fvQS���Wc"�
?��l��C�m��O8�K^%�� ���&�����e^���?9�R�5��'���8M�y�:8�qFM��h h�
�H_"_�&f�_H��0�{s�ӷg������e ��@������Ϟu�Ï����o�8���=��H�f\%����v6;Q^�Q�s����QP�\J�K�{2:(���/­Q�c�9�Pp�8C��Q�z./�J�G��G�:q�."=9�D�ȑ�D�����Zj��%��E�U�\�S	L�ô@j8�#�D Z�iV`�/�3
���� y~��뾫(ȓ�$�s���?�kg|�ه��#|SQ\"�g�y�֠h������Y�Ҫ����1B�($�ǟa�^r�H~�O��M:��ٵ��\$Y�Y�t&�|�܎H#$�(�4]~����c����ӧ��C�,tvP{G�Ҙ��ƑR�]*Z�FʄX���bɮb\� ��A�M����2|�-��G]�ET�8�� ,�P*u\�=s+?�kgO����l�]d�lX4	�8e���,��ތ�˩���FZ�ǱK�Z�$�afs:J�7����l/?��Lʍ��wh��$�L�ϓa+�ʩ���1÷��+Irm*���]�3Ϟ�EqH��s"g>��9��PI����1��&�3�f��sG�KJ�2�!��5eM���^�)�7;/r����(�]^����'�;f�W���'.������G��azp��� O�x#œP���CH
"�5z@��������%!.)\���].+BR��ڕ�J�<r�Qͮ��8����`��[���3�<���Η��o�'�������8�٠���-����D�������Kg�o��Ǵ4�r���F綖h���,�ͨw$nPU^��N}��/����w�;fx\����,g'O��ş��3�y����澊�׭��F_RX� ��u[s���La����3�=ꩪ��M��3��\0�S~�l���+7��߿��^;��Kg����׎�'N�zai����k�n<]������5��q:9�����W�{3m��Q�9�����#S�� 	����A�ɜ"��JNZ��|p�����_��ѓ;��q���ZZ*��'|ݤ��_����c������Vsi��    IEND�B`�PK   $d�X/�iz$  �$  /   images/2b96fa39-ee03-40f5-a6d5-dd88ef9bf1b1.png�Y�S��>8ܵx9�
o��ŭ?�݋�N��(��Ŋ�{qw-�?��L�ٝ�l6���$JME�  �*�Kk���=�u�p�U~�0��u� �ħ�u$�ݪ�W%���gwM'Kw/W��������������U։% �H� -��}���J23�oW-1����|e�D��6�d�$Q6p�|+az���m�';���nDс6���.ǳ	�2��Щ�H �H�3��f�|֜2�.�"��|"(���1�{�r�p���6.����Vp?ᦹޤ'\BAA!�4 ;��q�mhh(��� Z^Q�Z��!hW����㥧D�y+���g��29��8h�mL4D�f��z�p6�c�z��p�����=�h�F!X�T�~�YB�ԯ��\���{|�}�v�]�I��y.�_�p\�Ǜ�b:������ù1ا�����{��O�f�pwP����r�e�M<�������s�gX��Y���D��[�E��;߬���f�qW�`���=x���W�SU�|�Ӛ7��NmןƿK��VOX��^M��6UM�F�(���4��_��}|u�!��˾!�w'��Ȫ���n3&�w�(��K��Vv/c�*������C�s�n���f�u�֚=�n�����z}H���;�<���Y)þps�*��F����������W���z`�9N�=�����?\5�_�M��ᐃo��'f��ft� `���z}�a��4��ۺ���������Y� ���[cA��Țp|Z1��V�J��9��	P�u�8���*P����儲���$�' �{�i�]��1뻛3򭘱)��yM�^�n�ɞmDЮ����o�̀1�������jT�T����{�H�\���׃/���~T݃�k��r�{����=ƣL��H�Gn���ßq{�z���D Pë]ԩb��ǣ�`�v'A�kH��e�l��x]���'��I��Y��;���V��Jxs���[n�F�T� ��#$H�{�М���_�\r �j4��u��u�'Vs������v���ЖF��zΘ۠4���0��j�OnM���k��nm�� ������ˇe%�=
H~�:`�Զ�:BBK[��c�^�ւ�nؕ7�QA�`w�͑	�#�c�P���Z&!��~~~0��p�"�G��k��g������OQ9�N�y��}eDI'1G4,$��ܠ��ץ�����q��xW�%
"��➵ֻK
�/��x:�毵(Q�I�P�K�jyI�b���۠q|�a��?K�����%����;���b��O�s���N:����*��]�2>
�(�n�Y[����=����2p����$3t� ����U*o�Mn�� %f����~����R�u�����B�g�l�g��N�S�Y���ג<�
�GH�w���s����i��W<��^86��/�5�3\�1�Ժ��z��4��,Ӊn�6��DUx*t=������j���>����o�&v���U��/9��q
X���R�"�@^��O�b/��;b����rym4쫥���]䔬�=�1��Ɵ�.�H���¡]��`���w)'5~E�7��	,2#�ǥ���<�@��%p�(w�\�{���-�%�h�~�l�;9�h��� ����V���Z���x?����q�~/A-�L�>��OR]5���_)jm4�]�ۺ'���෮MI���T�o:�7c��!�ʀ���S�V�K���7��ry�=���<Ǽ�27�-(��������Ӝ����L^beӶ��{��Ũa(L#�Y{�GFs �vE ���Lъ������7�vA
�I����mذ�� �̓��|�`2�&e�B���*�V�!������oˍX�$��~�h��-2CG5+_�~q򅘷e��"I<L5�����)%�)�s$(�%�t��w�����J}�p�Gc�D`<y�co��v���h��k,G��y~QTω�`>ԟ��,��3�=�Śȅl����@3�!�=��Y?�'��K/�*~�.�;g�����k��7�c=����$��	 1]re9�q��q�_�MY��] ����Ȑi1��AT:0�_����}�����4�<DZ��r�AC�)�Wu�@��SI�^�\3E�"w!��x����J3�k����a���d�r���3jdL�lԿ�m�Y�:�a�<�i�f�4EE�DF����� �%�����QƜP���'N�5v%�Q�66A'��|)�)�-H���o�8�{�a�6�)h�������$��DfI��8$�g��{�e@ܬ���H�;c0<a��`~ի�f�^!�U�~%�>3�ߧ ں��N�	,r;\4Q��I�Y�W"�9H(�n�w��ka��l	��>����A1� T�� �QB#C�^���8���
����������i�Ꞛ^1&�t�;��
�ُ�iLK��;d��>� 6Q�C�y�Q�V���7�`����BXwW�қ$Q�}���Jۨ`��(8��p%Y����Q Qi��	���/��ڃj%H��2�M��<a�] �T�N��S0a�g�5�=E#؀�I'�r;�T\���\� �0���&�c�8:��Z�l��� �+�&?K��Rt3�/�|I��Fe��+*�����R-���Z)@Z�O	��4��m�S��Y�r<�\�B��fϲ��iF����; ֻ��v��G�B�q��3DK$�윉r��P��pI�m��,�������+�t1R�=���$p�-�Rm�#�B9 !�G2b$���>����Ciz�d2����$R �Qvaef�`���E���8g�	ˑ���;��=�p5�:6�������r��"�Ԍ��԰�$p�� Sz�5���(V����?�`�ƺ�ݱ�R�%�H�X ��@vM��Nfۏ�gX�X��I�l5��.Q�w��ㆵ��p OI���_x���o����Cx7������7e��{?�h����o���k����#�������w~��@��������4Fa��)t1���n8~"�4�#�uF���<(d��)��F����K�;<Qe�n)��$�X�
TD/���K���`���g���P��'04]	p�"ò�-Ob�6��+O���{���}�:r�K�6�p�e�� n`�鯍LPn�I*kRrx����ėe���<�Ĕ�P5L�q~AW�_�͉G�ߝ_a/Z�`с 2E�^�L6��HzDx��ľ/�\\�|���B{#	�!��G�/6)Qh¼����� 'A�.���ԧW�f&�;�E$�k�&|�;7s穽��Z���ވ�o��<ңc��v��M�L�i�T+�x4*Р� �:	0Iа�j`�R��Dʞ�	�
�/�z�^4��544�9F�uw�M�yd��
��^+�J���wg��]4\�`�ڤVR��D����PC�5�6��!'��ܯ�͂�����9�� ��*/���G�+�V����T-.H�Z��D!_�Ԥz�,�D��`9�����s��Hۨ��z��;]���ǟ�"�q���B�W�9��>A�NF+�j�/4�g��΍n;Ø��5GcB����;X.Te�D�ºc��[�S(���t*�~`S�:��D�<|��k���R�u� �����"#u�3]l:�J)؁\��x�<�<�ցq��3&�(���9T��+��xH�#F��u�
��U�CVɀ7�ش��}���H>V�k�1yL���o!J��	)'�ڹ��]f@�˹K�7+�$�a�{d���G��5F��NE��֑dA��5ߓ��!� �؍�i��r7R�˖J�:�\9��^
��T���~1�,�Ј���ٶC�~D��*Ƨ�������zs���Pk	�PG��G��냭MLRx)B�H�ZR�(�ӏ�:�D���YmI�eW:N�� 0y
��׊���6%�r�b�g5��o9�+��W��&f+I�l��2V�c0����q��ڒ��5q�ʏ��<�D��]��Tqx�14u�"B�z!���C��W�ؑ~��熹wj�|��O�AS�ЊC��2K�g����)Pt� 3s�?��@$��aRg�Τ�U"8P��+#�|]��o������t~�?w��vRy�*1��1�B�(��5Fy�D�Mn$I�}y��&.ϫ�3�%���Y��=������߰׫���41%�JS�z�+d���[�[&qc��ϧ����3vUC��O�$���W���
c��5pܢ2N��~�kl凓8y,67I@c��:V��hV)dH�,@[R,����Q�p��߆6��xo`TDU�2#����,f��D_C(��^�铅�� ���7bB�Iv:�Ͳ�_��.`^��|���s@r>yG��:\؆ ��j+�.����TۢN]*֥caQϵf|�.�f�\OQ�^:�IVZ���l����EY-��&�$��	�>ʨ�wK3}h��Y�;�z�4�(x*�D���rf	��?���nmۈ��3J�	�H 
D��ص2L��G����=��D�a��'���:���B�I��>�[�n�K��p3"u��Ͳ>�{a��H�
�ƚ�{oͰ�i���s�Z�9nfX;vN�Iۊ�������s6��d�����Ԗ;#ou��P�{��7n�ݪNѽJ��|���i�M��7�}�Q���>�+��m�9��,�Uɟ�69Yq]{��ryIO�^���_ȧ�7׮.�'��pob�1=H�<lF� ��Ȥ<�v1Z��_�}�^k�B�~�N�u/R�E����9��`&�~��\������u�z�����on:��L��T��G��~H`��u3C��$"]A84#^)Ջ��Ǽ~�<j� ���7��k5��b�L���w��5t�h��^Y�C���'�X-* ���U�k�Qd��">�.ռ:^�q�c)�*��G�P�1WD,ZN?~���#��4���������íۀ�fd��X�\�?��Bn�<k�>d��R���U�(��R��0�h4�"1؆p�ч��� gg+F�ye��9�7��#|�!�}:+?���$~ߟDu�����`���ijlϊ�)8�B�6�I�2,�m33Ց�yn�3�M�d�$�<�(��B��m)��˚���mx�<}�-�֒�������P�U���E?�b��PA�sN\/�yb�!,,�+����3&X?��s�Y�L~'F�|t��^�c'aP\���u];��*JX���n+_�J�谂��ɞ ��y����2O��yLfD���b��#��چߵ�rS��o,�ߋ2g3���� �w	�,#���.��nٲ��	������[&κ[:=���r�G`� �b�x�0B=d��!
ǵ,t�p��J�m��!|̆��h��N�]$M�֠rģ�T�.����Ӡʀ�H�Ǹ�5^�d���Ňm\�O%V�ͮ-:`��B�Xy	v����!��脏�>��"Ǣ��q�vLy9U."��}"���Ez~"���2ԽX��c^�^9&{�hs�V~�f���Dw�`AJ!lVD��Mx	�V��x�VX�/� ��ہ����m��;L�}r���r*5mE�_��B��ق�����
�&�z��Szt��u#L5/L�T==�1�:�>���Ȼj���A ���-�TH��k����䕒i@b�|UÚb[��Cʨw�_^r8IS]?Ԏ��	m�_E�z�=��X%׮p���>�yK������<v�����]Ѷ�G+��0_6�fi��v�DLg�m �����6�/i�χ��d��q$T����vg�g�������%�gn�6�s�_ː-fjw1"���W�ڐ�2�[N��5Fx2�dwb`�4���C46k�[�	����yk��`���5K�����~$3� 9H t���R�)Mt@Dy�G����N^�º�C�y�h���|�j�+��i[e$�,څ���(-U��ZL�c�K;m�2��t"�V-�)�.��SX��
e����HÛ䁄��)�䙱^�!�4/�T;�)hL�.�ܫͽQ��;��e��F<z!23t>���y/�:
qj���8�t{�ej��_�Vh�\ud���J'F�0�R~*�۷䐊��`�TD�Ve�%�s��ԣ�Ј�lvʅ������>��U٠�BlD9���L.��ڋ��N��^�@����c�MO�0yM��Z�˄�S�pև1C*����b`'��=+��}lc�|dr���I&��ekX�7>��_�|'�c��j� ��o';����K5KF�[u}����+�^��d$dd�C?gx5�R��O��� ��P��������$��W]Q,���21����R�=Ռ9,����Ed�����=�r�/�T����=��=�|�[�rX���x�P������a܇U�D:)Y�bQc+=���C�|�aҿ$���C�Y�WZ�J~XE����m�P����lm�>[_�j�r>��!�gɭ�}xO���˵)��6*�p�v���������תO��ьї!��e��$<��y`�PN��Q�7N]I���)��:c��_k?�F1�'<*���,���o�㱤D'�OC��d��}�2�&�As'�s�	�ED�؀!�,~���|�Y�i�w�eiX��>n��?o��׼<>H#��.`+����`Twk]�<)�v�:��{�|u��݃!�l��f�x�)/5x��'d����D�\e��&W��2ً�����E���#�����#ҵ:��|��_���;Yڕ�U���۹J��&7+�b}�:6Ad	6b���`��hNK=�)���H��D��W��鿙M��<���H��$!_��yB�;�s�����Q�v �A����ȹ�X�z�Q��������;䰪C|�)H��{t�@��;�\��V��*h��R!� >A�U'�r��Xon13d�s�޷b�`� E��L7_PZ�M1܄HMu"8�J����RJ�LY�
��i�yf�����9��9c���ҳ��gG������߇�P����π�� ��ߺ�9˻z�C�>h����H�����e�9�}�s�^���L�,�z��a(�;�`D@#m�D&�m)Z�$j��i��vbB��z�R�w׷�,/˦��`�&�i��"3�#x�"J�IW���56��u� �qp��k�S�.����)�vS��"�moe}� ���bG?mtd�-�~N���x6��j��',��f� �V�)�?��W)`{��ͣ�}�
R����DK��R���ڷ��0b�N�"em�#��������79���v��{���,��L-+��S�62�Ww�[�� /�c�����K-9�RUki&��opBR�'�a�o���Bη�i��\�|IG�F��DN[/��x�&Q^��`��������H���$e����d�_$�p���<�`�@�� J]\�c������N�7��	�����E"Ɉ1�
G���>Y�IV�ڷ�)e0*\����Yl5����=g��h��/�cRM�=%�Fh 9�eL�R�*u<�[JM&��T�i��<����
C�ml<����V�R�T�sDD�5kv���6��<&�w	���|�<�2ԇy�j����|t���P����_8���7��'�S��C���q|(_�/�:��Y�n��ׅ�[Ь� ��F'�ĉ��#!"K҉{�63͚�K>�����VD�2�Lq�S�����Y��r���?Ϯk�5��$-od@4cvP6�	��ܝmX���L[l�o�/K�-%���K���HK�*��ny��ޚ��n]�n����]Hib�;T����s'�<1���{�L�ҵˮ1v�h�C�g�Z�INُ��D��������>��w��E��'
�<]���4�a$�SP�q�
;TE�Q4f�é3lD������I� qü�~��g�57<�|��жt�4�d?��=��8G���W7~��%[y�g!r�*�g�:1��7&��}�+�j������	���f&�weO
�jYX�U���Lӝ��騂��^��I�V�.��P�p��0Jِ X�K名���@3�˲H��Q�R��Ǚ�XGT+���i�;��?��)�[�"��#~\q|0ϦY_l)�k���wN�B��?�;wqM��$����ƵNk-������������He�
���PA�P��h��a�2�,K[
�c)�k}�tɫ]������.�B"[��mp(<)|��������`���*���ӄmE2�V�U�K�� mL
7L���^��fԉp
���y�iP��+��j���H�r$HG�qq�Yq�~bbE�stM������ȟ�O�ػU�T�B���фK,(��%����d}�u�����aO]�N"TlԔǙQ��� ���)�<H�.�/%z0,�1��Z�ҭk�c��{1_0�.}�?��T��wzVW��EB $i����~����q= ��\�S�ݹ�2�j��l�K�B��g�mX�ۋj�(�-���F�>'�s��W~eg~�.)�����-�mQ��I�+�m�b���=�]nV��v*��S��9�ߕ��X���|�(�8��:��٣�����=�&��ꄜ�����$[*��&�[i3��bm��t���fxY�r%#���`�\�p�"a[4���D9�M?�T�^�������ݚ��,�b��p�(\�t�rf��+2��r�^��d�-Zw/���c<��u��/��I�h;�>�!���P�[�I�(���Z�B���ljj��h���7F�+)�#��%V��:���]�E^3�?�8�Ao|,&5Mm�Y	
���Ͼ�\\�3!j:>��2��S�$�&��m��6y�?�s�sJg2�m�v�\�����O=�I��������]4�U[�3�V��&�T���m���VA"1��[ </0=l��c���WD�Y�٥ '��X�s�)w�D��+9�
�Ж�֐f�|M�c�G�RLKy�wWM�H�3��Ϫ�Z��A� T�k	�P��T8��HN�oS��`�zNIc�<��6+ϛ��;�����k���d�(��Z��%lllBΦ��d�g{�8�*�s
ڝ�sg����.?U�iO��P\)�ܕ9��Й�T+��1{%��"��@z���dT�+%���PK   ��X��@� �S /   images/2c28e0dd-d0bf-4126-a9c2-80a014cb1784.png4{<����EfB�[V�2�����!{�l��;{DF�k�B�&��+;][\{��?����<������|=�����p�����(��,������ܺ���(�!x���?xO�w�o#��/�_#<�ݬ!����vN�pKsk^g7��M�;�]���3/����ߴn&�6< S�ng�"����R�;��QQ��*A��6.?6?.�.�2�+�o̑k���|z��b�R���^��fs��A�m ψ��k��ذu~�W'�sjX���,8	�}�����������	�U��D�X�voQ?xc<�-���6���h���	Mrļ���Ű#��j�l�%%�HXKJ�/��I�`kU0C�w��W��o:w�9��n��5�+�ᡋy�z:Z�t��%��C &2u��:>�zk��X"�Ou �w��Z�j� �.=z�/����ھ&G2�YD�F��?}y�n)y�C��*v^qH2���ffo+g�-���h	v0�+A�psۼj�X0L��ϑRS=S>|`z'w�S{!�1�7IJ(���g��Tq��k�@*�gee������x&3
��W��H)�.����2>�I��@�m��X��)u�u�����%����CΤ�U�1Ҧ0�����(�*]]]˞�	=]݃+Z��-�Z���,_�Sb�����{�����
��٧���5�Sj�C���1����t��J�4y�D!�ۻK��P���	�����:�ދ����f�D��>���=���X[/�u�moU6Q�%���}"f���	=���<r466��t+m������Q����s��`�H?��=W	Ǫ�����%(��������RQg����s�桺_Cy�����<�)M&q������!��*E�M�e�_߇4�ױ˒��>|(VJz�����jC-CD8M0+��<�4rS7�,p>][[�1���?�mf˦4&!�:�=0[�~,^�r'>#����v�S56VW�(++�T{q+��׈��ODHH7�q
��z$���3�}��Sydz�2!�Fk[i�}����*�恪(���H�T���<υ�v���NEd<��ZHil�k����-�P�D�JG�D6Χ$Z���XI9V��Wʻ���J#���Lt��:I�I��Tx[�wQ,S�NOO�����;2�cX��B5P���.Z��`��t��<ճ$Ol^��,a���.KB���3��
���Je��UrP^B�X�(~p�,���g���S+���<D��)��-�j藘�/��GN����`��"G��.4��ׄ�����%(�>�_��sG���zC&!���k[[�/9h_���L�zJR\��N5�d�̦���N��C������������-�� �kes3`�xg�I��y�avY��=ӕ��6V�F��l�㩔8�C,���LRL�iO�H����@�sȌ>�vww�Jiq���74Ĝ�����
(!�]�49t>���>:88�TA8�		yL�)JJ�;ڍ�r��珎�>Z�V&J���?���a(�,�
��P~0D���﷕U0l�z�{�pJ47-٭B��õ���Άm�ʠ:��p������>ݣ�� %�M��ᒳq�m��zIX+�SX��#��!A{��=~,=49ٌ/����u싁���7�߬Qt��Q����[ZZ,0�i��h�T<�$�i7Q�gUs<�.����u��S��6�$;��o7��a� �-��2i��<^���$|* �u]�S]UU%�����1.g�{3��MG+��s)�C�zx��
┆����J$��8��`��oví� yc�m�$�9~b�h����8�7p���Wׅ�
&�o�	��ԙ�͠kHy��{\��}9J0;�_�m�嵵R!�����kb�j��W�h.G�H��g6��k��,)���m�!�y`��?u�3�1>�L�s�a!˥_iYO��|7 �̾�<%���]@���B�R��i3���S�O�`(if���L ;��?'+0��̶+�w��R-%��*�J^���[�n��Ih&F3�i%8�m��[��.�c��8�w��)]Iz���4�@&m��ol���[F�Y�-� ��S�R�?�Sm���)��	*d�)Z�c�Ǩd.���"���5�J�5���dHh2I!�+��� r�!Ĕ��Z�8e{(H���I��+.��� tY���̠5f��� �� �)�2(),\"�QTG��{���ijdѯ���BA�W\Q!-i�F8MT-�@�o�{�|�T�Es$��E���t.Z\��]�nܸa����v�1I�lN5��z�*E��3  �[$ע��\��@$v4�!��d�m���eq�����]���e�YX�v��i!u&1�i���%�3�|E�+��Q�Ϡ���,{�A���j�:��k�=�Z�HYE%��]��
lJ��7��b+�xy9ù��)L���ͭ2���y�2���7�����&@#,��;�"��Cs�P��%~z���*:
��������==5nf�$��3\�v��v]:�s��_3'��Z0�6�u�{(�v��vd~,���?�-)���{����3�1e4�_���T���]:��XO&��<I����ږ4��p�BЗ�;�l�Z�ɉX��V�!������+ŗ����`3�φ�vQ|Wc4�;� ���=z��#[y$��r��9�/�zDe�݀u!�T����fZ�5tc�������ޚ��Vyb��ӳ�s��k[BF�E��p֩�R	���
�}��1�1QmR��?B4SRR����=/u���"|Bq�W\�U_8�~o�a���=OOO�#)�!.���:���R� 3�0�A�s�5�X�U�H�(��"��y����#	Q�9���\�^��6��k_qa���k&E�%��xnNf�/0�xi���A������˃:e�V���}-e5����ԑ�T �AT2��L��/kmm��U��k~tK�hg�}m� *(Xt���}B��.��eUҎgS��^#� �u5��nG�Sُq⃰}���ޠ�?�ˬ(��g�����vaO�IHԿ���vO�޹s�Q���䗍�^����%�q�p_������R&W���r�:^r�G5�$�8ɭ�n���~	pN@�?o��ƳH_��@��%O�%�rW4�f�+ěp�_�e,��r����K��v���1�pH�B/�����{���o��7���	�J�����_���v�io�u�a�{��/���R}0GX��B��*�h�k\Ei~~���sE�>@ʦd���BK_�IK
��������8���`���Be%�c����,�9|E�&�=��f?���˫��rC�$�	)|����KKQo��D222Ԇ��i��=�q<����gz���_����me·�͌[�||Qh�4ջ�؍�5k�+�/ �~1�|�F����9�������""�O�&�.����0:CYoF��g6��������g� �N���� �?�AV��)��4�*�6�\J��o/-�^��y~/a{���K�kt��ҕ)��}�4�����*���T�? s���}����] n�JУ���Sy%��ܬ;���Eq���쳅���Bsh+���=�Z�A�U͜��>�� w5!�N �D�ٔ"��:���n@�-���%%���r�R��y�\w4F��m�go
F��� �?��� �h����m.�S�d�<��Z��,:x�j��\7�^?�Q7c"p~�ȳ�}��t�ӝ��~��̒�*����&ǿ#����d��{���GH��Q������Z�E(���}{*��"�o��cf�X%�)����bnK�|1�V�}xyqv ��vc*���G�bv�?@�
�dA����$@�,�x��PĲ������UOz��g�7�t�}�g?n�i��^���{�A�r�k��5��s�8=pE1�Ϥ�WW�U�6s?T�-����r�ρ��(Z��z׊H4>�2��_[\�"E��$�e�Ԓ
�6���ؚ6��kbb2���6Ue��4h���󛻞�(�mQ���N�X� g%KJ�?��^�bE%sےc�
�H�0���A+~W��>��H����@�h���{&��׻�D��zJ������fWR��\T���"~S��zK��ߏ�җe2X�X�zN��5�Z@KC
M����{Q�hh5��#���[CɢGkm��~��%�Ѵ�V���zC��H^��@�紁���p�';5��=NB?���.A���A/`p���^4d�z�7��W�=n���*�<T�.*��x�^h7Q�xz�Ħ4�荅=td�}����L����Y26%-ի��( K�s�do���o�[F<��W���;�ԻZf�x>�u�0ͷ���4���#	��<�DĘ�Âd��O�;��¾*ͮǜ�gf0\�3{��q���!H�8%$����o;n�4�B%V�9 �~^^�L��]"�����'(��a=1G����[:���y� Hz����I���Rb�O�
��'e�h�?�v(�+%jp���*���'P�����מ���e�op�=��.cŝk�9d�b���L�����Q�Tc���>+}S���}?)Ӭ>�ri ��j_:y<g���4�5����=��3�Ȧe8��~|��\RR\R��̹�9t��)k]Lw��hl���-��z���k3<t1�8 �w�^��%��	�v�"��ie���(ɲ�c�Zc��7��	���Ub�u�7����DP����l�ΘC
e;��]X�9�t�]o(�X�Z_00c<�=�_��N�u&�44�ռ�Kaa�Շ,
�ڭjǌ_H�ׯ���/�v�]����*I2{��g�ًbQ0�� ��M\ 6.��8E��?:bⵔ�j�7M����p�P�8h���Z,)y��D�bK1��n��C���y�>L�����6�.x�����d��Z�C*�u�>����'G��TTPy3�K�gh2	�;F���w}||�ka��Y�я�˛�~𳸫��Hr��=(9Q��$��u��]̓{�~���̾�/^k������j����|��V�ze���e�3�V_d�V-3�d!�ر%�U@�w�䶽ٷ�8~k�猦��������[&�.����m�1��G �7fڮ"�uJ�t�,E9���B�~'��<u�Ԝ���h�l{0��C�<xPS�!=�y2mLw����1�e�?�O��p���Qa���^���o�� �v��W������I��`]��.�'�9_�������,����-�� T����.��:����&ӵ��/�FG�\4�����蚼x���&<��j{�k�f&�9w*
H���{O��ʏ��,�@��x��ۤ�X��T���^$����hx�������~�pj�A~��8���Θ����c�h���1G55�l�L������69p,�Ƥ�Z�u��w�e�Tn߃Q�@��ܠ=�NQJ�B9��~W}��#�ۺ3_��ܒ'M����:�Y��$��x.�,�bV��V�@Mkڊ�"�r)_�����3�H�K�lTz��0��\�pV�l���=�h8T����OO�RE�4����%�cY	 ����h}b�ŢJ�ItsbߧeW�?o;r]7��a`q�}Y��r�k�彴�K20ќ	�~��V#�v��TD��dm1*��0��H����M���Ԉ�x����ɧ��Ҋ�- �� -����+�YC�C6��u�\W�X��E���	��\�9|�,���٨g��^>kgy����5���F��bza���j�#߻��{�����-�rzz�A1����x���<��g���u3����=���� J���]WzR�U�ܼ/�\���c��s�]0.�ѥ�9�-Q �GrX�vN�M:��'-3Bl�I��&
<)�z���[�Z*@�/�]�I�E�K�N0HJ�F`e:`��'>�'@�R*'��ђ} ��r�q܊�� �@
�}��+��0V���߭�;��*NMN�s.���������(���
�q�w��t����m��m�yY0
+�v�̓���,����B:b��$�6����S�`�<~b<�W
�.>����yא��W5\�l�7����p��2�!��
�Y*�@��܉/��v����+N��,J���e7�,è/�c9�Ն�o<��2i��/,|n��,؞���
�e[KK�e Qo4,򦁶0Y�4Ո��B�2���/..�Sjf�����w��CU�E����t����Ө��X�	p�j9��LN6� �$<�����Ց��7쭻?�C�xr:���n�����'zK���1�G�K?4	�!f�ٰ�ci��OpX9�#E7 �s̀E�0�Ò���٥/5���|��xs/A�U�zP*�1�����
�ji���3g�z�s�s���(A���hV���*EА�{�r�E�=��}>�Mn��I�5�t�4h;"l����G�r�\o����;���� ��f&���l|0eK��Q,Ю��ߑ�.���SBj�ӆO���h�u]�>[wϊ��$�f�1�i@����?V�Z������dbb�  �&�m��E�!�9�bF{.C�_���M)���c�*E��>�P�ǡ�c����F���R�W�*��g�^���@�g9�A�������3�,	ўx��o����t�ò��=<^����q�KT�M`Wr�{&�cmm=��/i�u�
6�..*�V��eT���1�4s|3��Ŭ{��tL�f K8�1�@�p�n�kh�D��pQG�;�Df���PJn�m]�_f,���X�K[�n�+SDPJcc?�[R�:�� ֛kjF���E�*Q�����2SD(%=kU�"����؁�A��b��ْ�j�,�{;<�UP�h+L-\�:�|�6>��%a���;+�a\�C\��������a�����ё�ҦbPiҁR���a��zS����s6��7��˶ �wqk�#c|�nS=!�{�yZ<�gG��$�-=*=�}���s2�M�
�;���B��936�|P1N���{E---�`����0NMe0�(��eζ�GD]�^@"�Y�|�R�֭[�m�.f��m̜�<�Lp
*{�qv��A�$G��?�o��[me�\M9-�	7�jdjG4�R9�9gAb��v�~i�&A��W܂�'<���Χ-TM˛F��T��B��t�%;/��ZR8����z�� 5}IK{�Y<M�y@S̔�W��!訮6��iT��fD��ԫ~��Z +ilJ�0T�u�շ��y���@�ra'y�� ��{Wd��9�!�V�[\�P��v㔰���ן�Ǿ�����T�3<���Hd߫M��F��LoV���ES�~�a����XI�.F�w����w�Тe����H��X\�(9bNveN1��=$��N̰�8����u��G�ɈB�������?��s�.�y�ߎ�"s�S˿]����e���~�t���RR�v�Ix�fm`5^n�]��Õ��������N�i!��n)*��_f�KG��zO�=^{��L]�C&c�^H(�E��B�tS!;�`6��l�Z�s.��F.ތX�fk��m�illlMT}�0�Z�ԟA���f�y$f�
6��[/��p��'m�3����X!�ָ��PO��A�����ò�Ӄ5�(4�|N��}��?/q���C)s�F#א�:K�G��nuݵ2H��=1���3:�#�:-�I�mn���`�g�p�&� )�0Іʓ��WI��&�<���j�~*-E�X�����ϙ0��8�{������b���#(�NY_M]�}h��N�� �=e4ZK9�`=����v�mg��;�NE��F� ���Zj,Ƕ�����h5�]mg06�x8�z拍ɆR^۳NҞ�.s�O--"=�rG�0��@ ��g.��g=��
�s�%4���v�,h��?�<DK�N�IX�l
�59h_�
+��6jܒOPz.�����1��Z}Rs���@G[W�:6M= ����vܪz⊃��&��9�a�85(�����2^tru�?V`���7�v�C���pn	Byh�j�Hj O2ywyc���{M�a��|�2��QR����O��Q&�!�����Qʢ�i�}�DනN�G��/~R٣�O�>���(����In���2?<�&pI/3�S�@,�����C��d��?ONO�c=��7�:�VV��(;@�=&�Y��@u��L�kV?h�늨�A��eÞ��[@��re�Mb[y+�������s��������)��+B�bZ����y�����}���=��a����}K�6���n��sTWd�(ꋑ��)p�gG�`u4�ҲW���{������@���ճ�d�ŧ�QoHN�Ζ�m�KJ~���;u�|�6 bUI�Tn��U��ê">V���,�9Q�ƿ���I�(�ԙ<�^�ZG�>�.�ƳĢ��	r��o��c��0�Éq'��b�|��i�l����� s�F��'Z�� ]4�z����:r���I��[�]T.�(s��T���ڍU_"�!Z2y��J�X*)�)�Jp4�����"�2k�#+r�JT��l��#�=FO�׼-3�wTN^��j�Q���<M��C�����L��d�!����\`��B;�.�ݾ�<�t��8���2c�����*�56od�tD�7h����+��kA�� uz��Z�	PDupp�i�bX��e�W�l�~�|��!�`�\k��ު=Z[[-PIwK*jh�>�yǰ�7Z0�5 JG�%7X�KZ��#R�@�Q"e-��8{�^Ӣ�(Gm���4"D[��� �2��m@�Fq��������� v���*�ٸ�bm]��i4!5��ؗ�W+`�Z��Tt�`�7�˴9h?;y a� �+�yY'C'v��19�Rj�% �a�e�2#=7�<�ڀy��1h�a
�[xo]�J����=�q�{����,ۺ��4&��΃Cbm���$<�[�����Ռl�>ي���_���4Ќc����g'�-�:zz��|�b�7�g�|�ı����s��]^o���}'���\����>l����#�%o*�UJA�-�����ȽL����lP�P5�l56�$9,�WWwE��m���.�;�I��\v�$�В�s�+�{�Ғ�9%lk��<�&�����'�i`���0���^׌�]�pQ~�.�v��#��������\B���O���B��T��į�ۂ>{+����7����V�Ļ����6(7�u�1E���r�����r7��k�~B�7Њ�������VC�ԓT���H=�� 
�t�K�I/��tr�.JV����\q;��r�w�(s��a��C�2cW�L3P>ܼ
eee�K��"�+++�m�p�7�٢�y>���7mp�A���;ʃbf�r�zJ��n\)��N[D�Js�s~�ȱ�'j�=Q���`4�n�R)�-���k��M��)����G�]����?���M�ާ�+%��c�A#pDWjz�e�o�*o\-�%�aM���NNN�#(��Ps�\��'� �w�PDt�{���i����/�ɰ:C�k��+AXCT}`S���fd)�1�f�}�9���W �^�4��5~W�i\��~Ŗ�t��vf��������:Z�5��G������8.	O�7̀�M}�#��INtJ���fZd�u����f��2�*��!k
���q���Mu���B8j�1<���n}
�)wo?��)�#z��kXU�|4�Q�e������I�w��#�BE�{e&-]���b�'�B�\�|]��蚅���"�v����Ⅲ�7�L�n��~YT~d�_���zx��������7��Ҭ��O9��Vf;B(�V�R�҅�;����׃ëO�c��@ՔD�<,Q7�\][+;Xvػ����A��oY�p)l����븓c�Q���	3+�kz��/����w��:w�?�y͖�H�I�����+��&��Ʊ��\�YK"� �C����?m�m�YJ-���!��q�:��R/R�����Q�x߁LS�`mp��@B�� �����pN^>����'~R((\-A}��L`�;v���D�����>�}G�9�I���T��) �ə�e_;�6�LKZ�\�`��#3��u�ra���M~�$����!S��F@��ʻ���x����j9�*Ql�&��m˔eX���(w� (�Y&I���<"��95�n���w�T��bŔ��������n|]�U.s2
��������ˌ���PqUIf��!�x�0D�x
�_��lj޹B�X����'Jɶ��l]T�t�"��H4�K������������-�����#�T���m�����xf8ޜ�j;����^Wɚ��4U�)Y����b�#Q<eX`�p��H���� ���Z���>QN�o~k�aC��|�z�h�xg��5p�yp����Yaa�,�j\�W��Gm�����ڍoFK���1?��W`���$���F6���,��<��{k�g��;���c�;A�S�r5���_��3g?��Y:�	�5k (���*�3��@�徱����M�1Q��������Zy�PyU�v�jI)cu�Uz�ߡ�*%��~ט�%(����� ���������߇���q�[�g�r�0�ҟ��IA$W��<�1��F7�t�������o�8�����J����|..v�E�D�K��A�<ۻ���Ƚ�P*�[��U%���V/3���b��c�@����8���5C���8�ĉl(���8�&]��W5otE)�^��44,5
8Y��Ht_�ǝi��i+]w��gc�#��А���,u���\p�%
 $.��p����g{���6+Z��.�@&r�!A(�"%%%�*j+�WV�@]i2J�y���>"3>�+�B��]�M���7r�M�nb���$����8�9�7�O,��Xw`-���=>rĘ��=������"�!��V4)Cr�#����w9�mU���b�t�3��:��ÿKKK�L��UU�v}��q��B9�L��d#(@�ɻG�L�����}����vg����ʸ���w���lP,\9�Zx0�D6���7�k�������s�<��W�Qu�eg(��^O�ހ���y�q��#g��h�.�ڰ���l�D3��n��Ʊ���Z�����R<O�c�?�����X"ދb)�)t���].G���I�,Yڥ7�7�(3��1���@��͌�"|f������?LD�j� b�ym��6���R@�� �9Z#��/;�����'�R��߿�����|�h;����HP������j�X�#6��H[+t_d=��$y��ڍ�Zq�a]]�GQX�x�vq ���7��kr��aE�A�����2袃������c@�1=~@#?66��{�i�]l�I3�K��k+(�^<������)��/#[R2�Vd�N�=T��e�B�>��Q6ꄩm�gw�HR�]�L�]f�K�G��･E9<Qk,:��c��=��Lz�y�W{�ˣߣƼ&Reg��F�".kk�Ξ~R�u�NM9zzz�xMz��*����m�7^�)��ST�����e�V]����
P���(%Z������iM�X-�~��8ʷ?�`�)�ɞ�!��W�⿣�rwj+���`�.s���i]�}�3,N�J���:O��͎H���x�F�W]�(moo�h�oOm� Մk�oM��I��TT�<�?�O�]���~�Cڋ%b~�?�����eS� ���v�Pr8:��S2���U%��}�AU���\��D���e�����yg���������p�A	맂�Egy��w���ގ>C6�^�Nf���R��p��Bg�:R��7t۲��n|sy�kcS������6���Q�����h��|cH�z�r}VJ�������D�9M�9���Xh���w��qF(��*3ID)k�M�kfS��[�hp n�(sW'�,�ko�0}��N| L�#���?��v[$�S�6UW�nn�.��[c�ĤL�Am�4������E����r���NR
8�LW�%����DY&ס����+�&�ٔ��V��f�P^Z�8�3G���(9?�]�a��@<dSe��߾����ԧ�)���gȫ_��&��M������z�����^�L�x��7[��W� y���0F
�o�����0T�ތ/�!����z�zsHQ����-�}tsD0�����_��,,��G�GK^uP���ov�A!��a��)|��n�����2�<�t���a�P���6Ye�::䍶��^0�����u�>�L�3�gX��Y�C�3�	V�;��Vf
T���x��d��8�7����s<��:v�G���~�G>B7X���B�V#i���2��Rpwm�Žw�ݶ�cF-�J�1���y��#�K�|�#��1�?bepn����O�L�����T۹����-��XЫD Wb�M�s�ǎ����.���2�n�9�1�c���ISY��B�`/.�����40�� Q�r�im9�ח �jƯ���`�����;^f�3 ����s�'��RK�{#ޏY�6��
&j%�Y�8bZ�q{	�CB7�qDSk�v�9wt�E$�\ϛE>�Ԫu�rc��j0�}�AKVhwǉ�a��N�~~�s�:�ط���3�EN�1�F�9�<�����a][�Jc�v�b����hؼ_�:R�r6A��h��A���������)���lCО�&�o�;̮�h�4�{>:���XO�k�^�]\\��������yAm��_����b�̀�y����	;)`Y�Dֺ���#�����hY�2�a.�5L��v����g'J�>�įEZB�X%&l6�n�~R����f�+��H*����y]�?�X��-�A��Q)��=o���S�M����<A1FÃb����NҐ�Rפ* B�=O�n�F �s�n���2�M	(�t������D�C�GL��t?ct#���B���(5ӵ��Q4W��p8�D�j�ۨ]����?�{��3�A�}��oaa=WDЉ>^ω�
*Hj�up���Ȝ�:��y�_��wx��Շѩ�� idH*��p羅�]S)//�ȃ#o$Ì����tAc��ְ�B$���_��DC������ҩ�Sls�T&J#ț��~�N9P�ʐ 鎘8�Cկ����" [*���b�����.H��_��[Y�Ki���������/~�g<6��aI�_�m�b�6:D|�Ѧ�#�ע��r�L�D���`Y̡qޣ�:��5SJP#e���~rW|w�zF#�}u���x�K��料���޸t4�����s���P���6��S�<vVR�:~`@����Nt/� mԙͥ55�F媈��4�𗺺�1�9�b����EU5��5����	���%dH.?ó�6��9#�i�^�UxN��j߈7U@m�6��}�r���9���.�"RK�]6���p1O����mX A�[�J(���|z .ww�>�lV�|��F�N8��mL�6@"�z9��F}��F��}��n���)/������A���NG+��-c	��LLLqƿ��.���i�&1}[t��D�9��j�X��A'b�W�T������K#�9+���`�'vqL�%�~=Cu�_�����|�`p��b��E2��Ca7���5�,�M_��/b�?�b�ib���c!�+���������$nj����w���D�#&/r��Ľ�zC��l�����'��yxʜȶ�v+�w	����Cڇ��#o�i����Z��b �3�A��|�/����J��k\\��MPG�S�'iI�Tا��d6�H`J��q
�o���DϢ@����2֫P:�'��ͩ��&ϭ10D&��_( �c ���>�(���&�[��� R�7\�|LC-�����~����(��4���v��Y1���;;�o��J���qQ���]"W�[ S+�!�5���.���7���@&����&��)6q���r���n�`����gM���1�_�`jȥ���Y͠-�AN�,�P��k2?�ˑ�O�,�SXԒ����+59f��"�N��h^f�u�����h�"���9������k�L���O*0f�q;U3'��r=		W(O�\ϲσ�^�%�������n�*�E�2լI���?�h�	n�����y��U���Ԍ�m6`5�� �p��
S�#V��A�#d�|=��3��b�
�A���v#C�rݻ�"Hޕ3x$�Ayb��c�6�K���!w����m�a�-r�gg6�b�Q��|/EL�,h<d܄!�{,��925��#l����l�z2��[�v���'w�$E��u8��6���p�V����cP��]��l�x�q�3�耂1���t��9���߯���R���櫔�����Ū	��s<�(�0'�g�&��s��$������bݶ��/J�¯�2����rO;{�&�q�ޚT������q�Զ���'���V=�+�P�d&A ;�'=���.y��gl߁Z�0�]�"�֬��P͖2�&ӊ4ݘn1�v�G��W�ʛ�][�ule|��N��y�6�,gA���:�bc9���m�����ə>�g`�Lf�C8	3n�{�"R���4
q�H���y ��{�/`�	]���Pe"�,~���F�6n�^��<��)��u^��?�w<�ֈ�7+��[��h����8F�&�.�i�b�c`���L~�� �+��8���,��e 7ا,ا�篴G���� `��7Głb
�WTD���u.��W�b+G��?��}w�?0^똯��h�Ŋ^�ML���ܒg.Tۛ~�ܼ>=8�oa~�ȶI�������2ر��vP�(�.�Eo����.�{Pbv�>==�6j��w]H���H-8�Ro]OϺ�#'X$������m᩼��A���+�[�Z�Uˌ���h�0|t;^=���㦋���s������F����t�Nޝ ����8��1�b�h������j��^!0���U��Q��	�~��hyKK^�LIE��h�q��Q �Њ����M�����3 �Oqo됰&�ĦTC���Q�D��2��!�b��l��A�P�5�:%&��G���*��|�@�Kz�CM��s �E<;4sL�v�K�0�B���	O�g��uVT%��g�P����ҵ�X��~c`a73Ps����X���!�?٨�=6'W����N����#�^ӥ�~�tM��<v"L��B9�^����
h!�Iц����Iz��5��_�����y�t���6�k ,/H��t�`L%]��k�k�Y�Cg'ł"��>�P7�&���U��gg�6�`�ߕD��i�K�o����6���ټGq+%BgZ�bi�e3ߡ�>���"n\��d�L�Q�L�X���zz��^㞕�q܂SO�zk�(%��P�5(�����pH�\]���تrĸ�P���]y��:/�Nul�[c3�����K�⃤@�@A�MO,49&j7&�d�JZ�3�Yp�:����r�M&�}�yF���Ǘ������'\��w�:645��p������D��4��@m�O@�1��+^3R��ŀ(so�)����g�G�h��P_Sߍ�<��eG��+�(}*��.���IDNNG����Bk[�{��?<@">b�8�1' 	*om5!��b�}Q�������&�H6=��Ţ���a��fwpw�=�
1C�����fyk�sR]�j�S�9^n\�h�Z����ϑ�e���w�εe~��zʮ�����{����X{���������:��&Y[��'�@|^�3�ŉ!�R=Ѝ��&��&��.^�*b�:��J{���!'��\��誗E�Pq�y�@ܫ��ee�]|%OSc�d!A�`2=�+#�;�xh!�߬����������eA����>[���q��ʌ�ϣ4�ya��p9��� ���A�Z��lJY�g��cW����;~�y"SY5�^Rn2���+�m..&m�B�Ƈ�_\�P��a�h�e��;���4{�QQW�gQ��(O���)rzz�[�F�X��ptt0��b@	���B�����U""<�2H9p��q��ŏh���uF�{���ْ�Z�~Oo�t�>0FA\��-F��g�Rr�l<ԙs���6��f���SQ���w������||�W���^�CF	k�������O�ñ
e��%%T����X��7 �#) �GGmK+㴕WWW%�s��[�/@�F��k��ƭ�	Z��
�� ;�;B}7��Gߚ�C:�8ql��j������a��^$w����c^�%�8	؀�����_�z{��dr�͜C$k�CU�m��n�AΣ��cА���"��e�~�E���
��lS h���lӀ�<�lQ��@>9Z�f�"�
����c�,��\�~��mjj�	b�!�gs}�Aľ8@�A{��W�Bh��C�#d��'���	8D4i����k�vxn�k4���v�zaw-���.zlqޣcR����ޅT74��2S11����n�����������xi-�n��Ԗ�,R~�L{�g �F[��F��Y�}o���[��K)&ޫ(�F�}���+� o���`�s����/(:������sƔˍq�Zo�/$�<F�ª`�4�|�vG�"k�����lme�w��2�$�=�l=��],��A��ip 3r/���@�,�n��j�������f��Q𩰰'i��AR%���v�|!���P<�4�t[T��T�R@��	S�\я���rmcc����Ma#
b�lB�Uaz����@n[[ ��`S��#I��cPU0�� .�ho1���{�oL�z��d98c�{��rZ� h�f�2RL��,*tD��hq��:K����*������`Z؞�a����&��-��u/��%`.
���?�66~�9	ąP���`Zl�&��������'�	�~"m�1 ������Ǒ����b=� !s�x-u;�6x[���7Аc��Ώ]��9e �cobF�>zj��������3S�Ɲ�v��8�,D����4���{�@��a�� �W�Mm	ĭ��ɓ'4bظ��ޗ�CՇ�Ad�B��&Ki!����ۘB�udi0�'Yƚ$��U�,�}�dJk��Sa�-��3������^�^ݷs��s-��}��q�:��iN�B�L,���VW��e�ya2��n/ 1�Ng��������ӀdK��j�ٳac�F�U@nV1����ߪ��`��.��/�g�G+p[t~:�Qw����l������d���~�A5���t@����j�/^h]#���rA��x�I�V�hh��[�P\���.�2�/�vg0]j}e����q&�j�����"����!,�P@Ό�z�tarQC�a:�=����}����qz��������O۝|��,�
�#�H k�/t�M��P��i�i=�8�S�V����@�Mc
��2r�:5��ps_+����5H3��A�n$��z?�汣��/\�<tkn�
WS�,F�?��:�W��7��m�BC�Y�P�*�(v���I$K�}�;��}�h�rX�?�|SO2o��y���17�O|xD#Є�le�Y��p3��<�t^Ŵ3�us~pm���ş[VO�ԭ�"l��/���Wn��u=|1�Q�IpL�iֲ#\2��^ޮԺ�}�G}����nz���P*�m��ķ0��2����1&���sn�f"�S���	Ց_�hR&�4^L/���� �
z�=9�IY��R]M-�Hb���w�&��J���1y|��[-�1�٥d�	�}D/�"ju�h���dW�n3<|"x�pO^Ҍ��Z/%�s�2Ĉ=��,�w+�y �lB_���y����/��-&T*���pa#OkR<eR�}�������~OЄ�R��b����n��QwQ6�#G0啋��L���|ͨ��h�~)9����{t�����=�G��8+"�N�CB��_Hv��Y���ewvv�����V�Ld��zO+�%%����^}P��d���� �'L����V57�����+����V����1����2��*۽����Ѓ~��x��KJ�2��i�^�ij���}�V��R�JK��t����s�Ul(^�t��:��)�Þ���^$�����B����L7Z ��E�wOYZD�(�IX'�J��_�6�jX�;�Z���S]�.=� Ǽ|���_��$;��K깽Qt�Hp��t8HP���� �m� ;�A�F2�g���&!ߨ?�U>� TJ��$�F*v�3�'��Z]O%�A�t��o'�~{�lm�?'�/cʔ�Y���i�-���nŎe"��ѿ��9X�1HP��q�����@�%�ꍥ����I훀��F���#�ã���'�m`�H� ;G��������Ж���m���^�����r�C���WML�L��}^�M�?�Q�rZ�U/�b+t�d�X	�d��ࣺ�j�Zv/��H�-�s�Y�Z�U���=W¨[t(&��yz�m.�1�b8��|Y����8�y�L����n���sm�����`�+�x([s�|r�~A��?�#_�JӬ�Lt(�=Y�~�����Qd";�� ��~Z��h�.lV��[HΗ/WPb�e�7N��ESX���66�� �2�jcO��#�ד�����W��A��d�x:p/ ;v���Y��%NJ��|�ӝQ%y�M���}����q��w"��� ��Q�c�7.$�/ߔ�0VpJ���Wk�q���͎��A�����a�P�S��>�}�gm���Y_�\cB&�����o�>�P���<	.r�:�� ��_n�w�0�rr"��ON�?]�x�&�{8N	>���������4
&�TE�3���OʞV
(�X^&69C�MU�t�i=Ȣ���P���/�(5�����*&��g<S�?�m����8;ZM3Sx��/%�M��Þg����j:����%�w����(�=�BW��˪�/%c�['����[Ev�wS&�XO�ߢ�d�ç�v,�X�)��UL�����/�rj�Ro�=K">��ܡ�Zc��zLN~*dbM���$��G%{��|�r�s��q�A`�� jCK?C�U Q�����>�u0U(���
�nP1Eu���2
^\\sg����O��pX��t5�Q���(�M\�J4�����\UW��4<��j׺1]�Q�M�+rZJ��eMT�)A��� ��l�Q�Y��AN��A&��Q��gF��+߹s����A~�s\����b+ܿ:�~�c���R��_Lܢ���Ե��-��$\q�U��k���5��)���M^�n����S%3-K��	_#/��5|�KT���NO���::���Y(�/�?8�uP�x_&�d	O��/t�q�ݡ���LI��M��B�P�϶�t�d�~�(��2x@�K�hh��1��i�G�E�@^�o6�S�K���pB%z�Ӝ��A�_i���Xj�[(�ۨz�\��Ր���$:Gd�O�ؚ�����O�;���+�0;i�r�����$�vr������?���_^�ǭ�~Y�q�_]I����*��� �;���b:���~�H���i��������Q��X:uxY���mG1(�&�re]]� c�Z��vLV1�`���-K0�ݙk�;���@5��Y�#"��Q�T�P��>/�!ך�I��S/d�Wp4f�L�P?9ZA��5�߿Och��I2Ws'��}�ry�A�ز�\���^<`��]�|�����Ѐ���_��#��Qz�.�a�6	����Տo
o���iTO�n��(�ϣ1>X�W5��q�!��6x��R��|.5uuܵ�W��Z�E)��֗Է7�w6x��AP��of�,����ҿ�=�����T���3�lI������o`�!{ڦ�f��)NM���9H�B�u[fhuM�H��o����-�#��"4�^�,�9�=�q��".T�<'����F+e��dee�����F7,ѻF]UD�D>d�mOaʛ�i��� [�*K��س�j}�%�QT�M�� .�f>��Z�����_�(s���l�/�V��GZz\w�_oqB�^	��w[��0;%�j���#�"g�Y[������t���z����i�	�[������W�`	�f.C��kr���E1�7OԻ���5ʌ�R9�_��>'����L����42�C/��/���@y�ț���ܷy8�X�;Q��[8��`
L���j2|Fy�*�z�WO���D��-�5�qJ��-7g��b�S|�(���*���>��jp>��u}�&����A*���l

�@Ѧ�����/8+?Uݜ�l��,l��]O�v����R"G	����by������������@Q~S��6wy���?9i��Q�>_���D����K�Hd淌s��( �/_�<��NJ�a�3�--�Yf3��:l��%�5|p�����ᆃ0�+Eo�����w���k����8Qc�G�d���E��m�M�6�D
t٬��iG�eY��m^��T����l
����pc���wf�g��qH�����̒��oP*�{T#�m6�f�������ԗ��
��TF5�=��0����lbʢ��C^�y
��n���Y�-U�f�k���E��@��(!�����En^{%)�Ȧ/��=dny�k��j���6@&���묌m0��-aoq���p�Z9G�ꦦ��P���E�TD�Lo�@@��:voy�*�ư���eq߁k�ƚ�]8A��Ss�i_;ش�]Ա���`B) f��X��W:�#�us�Iw�����I�ɐ����V���>��K��'En�W��c���P�F݋� tb�_�H�2	ZwϠ��L���E�o,��¯?�5�\8oa���?)$���2	srr�E�A�v��s�R�׬�g���ֶI���F�R�sj^Φ������K�L������;�a~Ή��Dpپ��Z1��崟,��/�jS>>��Y+h��öe��
Q�ȜNg�Y��������bzL/z���t~��� ,y��<����ĺ�{�+��%R�� �?+�ߨ�Q���nz�9�M��R-�%=7��ܶ�	�F����]G�o� 1�4�vo�����U�����H�i�[�F�7�h�f]��LZO�Пdc�۝���vNM�y3o�2�+Â�N������w��0���Q7��Նa3�п�,��x5�Дd!^Q�>S�F�[w��_��ɶ�ϩ�7�P�l8IR�y���y�:�pr�DJ��UՏ^r��z,S�0tO���J}�lλ7��~��M�aıX�gyp�'�+��M���&m�[��@���B�g���'��"ϴw�j;�о(�X�[���v��k��8���l$n���|�ić�8�l��X��?<�rx[��@��=8=���C(0E�������ޭ�1�\P�?:h���zἺZn��*wn���0[���?pJě�Z�v ���7����d֏8�;쫙e�ȏ�����*暎̋/�AY�� �u˛��q��`|����L.i��X��x���ʹ���A���p��C� ��߾!@�<�i��:'d:A��݇kY2����E���n�V��Ug�|��j^�����?��������|�����ȝ7����_C��ӕ�>��ϑ]KZ���~�&t �wX�7���ɯg@����f
�O���!Dn�nU��B���A �в�8�!����z 8��;��<f&�}�J�L>�F�Gp�C^j��R�B��F/�]��C�%G�rvL���^�u�f���W��+g �{R �T��=��J$+�O ������	�b3 ߜ�h�~m�R�k�f�Y�Z0W�.�f�=�(�\��ax}aa��>=��Z�}Ҿ98�^3�*n!3�i8�Dd����n�Uꁰ늁I�MW��F�xCZ�����}ǽkղ�lT�������\�3�v:W���� �����F��R1��#m`�P�<{hQ�"��F�]���Rb걺
 ��� ʶ �mj��� d�/��]�΂��8�	��=P�0  c����g`s@0} [�A_�`�����s�I$@.�Y��'����1Dk�AF"Ѡgi��\�p4ٵ����A��Iָ�&�a�7��5L�(����E��R�����8��K
���X�bF�0�y_��(���}#��0O}��0z����F�H����W�#���/���d�	� ���}ŉ�}�B���g5� F���N� r>�5pF�ʋgkMB��z�t8�8R���҅��z��#~&($c�뱘;Z-�V�ɠ6σ}C[Fwy�N�Z����g��ρ�{��F��,Ɲkmu�Kbm���$����yP�� $����/Md�E�wI�h�x'
�O�D���Sm��TL��^��Ec$]1�u�(�v��SvZ��ݸ�����?o�C<p:7��>��Pؿ�ޱ��V�=B"_�3�D\����	N^�ܤ��s���5�,ʁ�o¯�K��
�qJ�;-Mb�#I�y�|<��ր�@���Z�A������_�574 �|%	 ��;��U3x��f��2�㚭�c����v��2.�[n��#Jq����9�����\��[ogg����u��-W�-f��&#��r�D�\Ҫ������� "}wEw;��UP-�<kY�{��G�`��+6O�^M�Fҫ�e�Hw~�ܥ>Ǎ��º2cP��Y�%��Y~sp��ΫF�J#�(�ɥ�&�ƃ���q�O�l>�Du�|n�E��P�]8���e�� �(J���ݣy���f|�}��.��}��C�i�W�^'��@�b�'��K8�����|�gG����L&_���dѾ#�s��IVz)��C��|s�]�����R-A�|���&`f%���={�I�Z?YOC��m5���1A�,^��k�J�d��<��S����~�B��L≿0٭}k�3��L`��4��#����TDP�@����bj�'��@��kv+��h|o'��߸�P8E��.־f�t�M�]�����>�/�>S���g��/
^��ȫ.�&$�׳����75�M����bf����������,L�,��߯y�/¬A�(y�Q1�#���lj�b+\��|��߫F>�tΜ�A�WA�6Lv�Q�	9�O�,�jh������R��f�n��<7��x���j֬�Id7�/�L���p���w8_ ��r�
����f!��Kt.P��T������DANM�� �����K���*Z�޽����N>j*����\]�V ��*���p в��0�aB��xQ�_�x%�l�l�AT��uV> ����ߥ��Y*eRɏ�w�O���r�)Ȳ �..Q���3���7���+��GgL
x�������� O�7�Y�f�,M�;~7�jf�@/<+��mh/XN -���J~w&k+��/����Y�L ��pL�кش���qw����S3�V!p(н�
�q��?k���|����dbg7V~5)~��=��|�|�܍��?`���f{�K:�J�~� �*s��?�b
�BfzVw?Vp��2�6Lຘܖy6�y̋t�Zٍ���@���>���i���b7�ܜ/h�co�e1y��^��S�A(8�ŹG9�B*~]S� F�����3���r�SF�'�lM�i9G�!Ci�B�҅>A3��Ϭ�wA�.\-�_��Ȗk�h�Aa��S��l�2������~"Y���8^�<Y�2c�h���P!��"�@Q���B�w��Q�T�ư�$σ��y������ܮ�U��ٌ���4����j�d���=H���A0w��%�Y�p���6��{޿j�� ��]E�&�LM��d�ʁ�s�u���{ۅ��b1\t0ϩD�<��㨙����ځ݄�$ɳ
T��V���/vE�t�B�~Cżw�$ll/���B�	�7�9ՈIt�i PX .�y�}nOŠ���D���-\���+Z{�ps�.�5`�\��*�S�נ��Q��0��D �g�"��뱒���Z�*��;��V��8��!q] WW�U���_��A��Q�|,$���.qn���M�ۄ���Fv�������f�ފs�:�!�X~&�|7����x��ƿ���Ӌe�<�L��K�G�=�����ƞt~R��I��F�j����UIKge��f�=���uD
�ޕ���!;s��ȅ��ѠW�����Ye�ʅ1w�	��+�� \��5�[�� r�5�#?]��?�@o^�pS(���z1�A߈�����"��*�V59���˾ɞq6A�?��ȀN��}/����)38;m��"�/���u�	1��@Ԍr�Ŀ?��"��lhg��hm����8<LGuKo�N�s��'ͦX3I��l�O��Civ�@9$�6���@���Pp�K����?w�9Ժ�Z<@Honm�>�ꕵ���աC��t�+n�t���tm����Yib"}� �pV�������;��)V��C�Woݺ=2lKF�P�m�I4�S-���ܛ}^�}�amaN����D��JE�����z����� �m��Hqp�ߤ}�u���-3��Z��| �YD"ߴ���)5r!����u:_2��N�9h�3��=�V��M��	�x��"�S���AeWL�ő�8�MInáȻT�va�v�R�J��@���(E3&���LζB��⾏�l�,�����%ȍDƖ�$��p�8~��QJ4BJ����3���Ъos`��n���Ň2@d�-A�9����ç߂�Q1E��%*~�|�ϟy��ʥS�'t��8�^�+.�d���q%˨۩�� ���r�*k�&ӌ1[C/˛�g�B���i�R�T�* ��j>������6&�v�ڳ��{ZS%H.û��v�r/���h���S���/#�\��Df��^�t�ףC���9	��>�d���싒�>|0M*8���{�R�4�Zrs'��y�p��LN=�yHi�N��bֹ��f �t�}�s���iHC���L�R�w��p���&
�����足���y��/VWr��oU2��χ/��Q�4uL�o�������vy0�~G/���!�����VcS÷0����֐-KH�1CW��7�$4!xR�*�\I��DK�wH��B�IZ��g�>�*�3��޵_k��Xg\�qa򣇚@P�iH�K�ۍ�/��!�J��_fo�z���H�a�y�����w���L+cRi�W2Yu)��}���¨� Y�gV�S�=姗���KSݏ�߾�=[��bm��k��<d�R�d�E"1(�Ї~�u�$ݹmC3N�=�L�y�{�TӲzN��c����*��W�n���f�)k��J�Z\��P�u�Yg-q�����V�,����8I��������ö�[�>������jO=Ş�,=��
i$ku���O�)�W�iǉ&zeg�1d�|H�N���PX��<t<��ٝ�_�)���7.�4������F���ocF}t�:K2Є���4�4�j�VZ6�Az�
���M/���������R���*��d
MS�=:�Kk#N�pVl�T����;��Z&���?~@9�x^�"_)�AC[r���0E��L6��!�ߓ3�`�YSb�H~d��M��'aT����f� ^�����m1[9�ǂ<k���$�5Bއ*��o{.����Y�:�1=��o���}��3�'/$�]U6j�E{�
_�|~]�xs�E�GW�ַ���^;�^;b�>�FX~�S���s��DC�u�U��� ���������ay�D�~�x����mcէ&�ͫd��W��O.��\�>��+?&�/,a�������A��c%&��>^�E�����S�Ny�d�4�2���	W$�x��ّ�P��9��Z7�?x�jȺ�mE�2�����塋����������G��Z�\
=�R��U4f�Cm�o���z5����yHQ2�:!(�v@Q;�|0�_|����!�;*M�-��(�-��C!����H:P$��Ӭ�?���.����
]��7��V��V>7�[�(�}+#�3s��%�}$r��$x4&�uuಊ�z�b�N'H�~��iz&��d� ��S .��utsd-�'*�uU��ˎ7�\��e��l>kY�C(�ds���yW� ]I�}�y�acH�ԋ��8N�Kv!5k����!.�2�.����=��¢�[��4��]W�@���
~AG�
Ɍ�"ъu�܄���ٚt��%-Ä!�!�&�G��˦0;BL1�FE(��B�}Z�C������;3�.�)$�Q7�)��6�]���V�uy�9�B��aT�<4[��������L�n�]��(��;�w�����혳����xڑD��p�������ֆav�B%�"u�3�G��CN��S��%L��c��%�hh���᩟�y��A�6�����{�.|n�^���gD_ن�2�"���=jH��ԋV��{�x�yQ��w���q��C�Iw^�B�I����Z�X��Ʉ�/�,x�%٧B�)���Ǻ:���7�y�N��C%�(��u�=��Ph�vt�;4f��\�f�S�A�y�������%����Ȱ��I�S��s`7���~t�ǭv���e$9�����U��= ̟���������B!�7�Q%.����W�4�u'|>7��=Fzl�N����N`������B���	���/_�jZ��=dۊ�1f�5�Ǎgn^U��>����
zб�]��g���<�� 臇��n�>��	�hfZ�уҼB��i+��j�7�����U����<��	����^PZK����� �;鋯�։Q��7S/*��B|�}RΪK��٭�2��Rz:ZwH-%8�\��3�Ҳ|���?���%�� ��ͦm��VƶM����������)��PH� �MO������ۼ��ǉ֞*�ރ?�n� +[�N�i^Y�H��ܐB�����~1Hꨜ;�<���F2�c�z;S��ǍV 9/3����X|:J��聙�93Ҋ�:�;dp��y��DgagW�w���x���*'X��F}�۰5�<^��|�2��mm�v K���{�,3������穜?bQ^�i��¹�����kU��N��$�����V�=��I���3���Bx�n��R�y��P�ҍ�'�i^�*��ă=�����eF�Z�N3C8XFO�hXY�s">�5ơs�Љ�<k����)�c���y�f����$�D���3Չh2͓��~��N>C��YA=
*��{�A�Ba���k͎��mAS��M�0bY��L\���
TXMK�YC@Da�v����y� u{��eׅmN$J@ �cײ�����/L0�[P�d����ᅅ����Y�%��S�i�k���S�� �*����wH����g^��f���m^���y<^<�-ɬ�lԟ��gB����,7�{�3,��64�@�:�+?���H,�E��%���B~ ���^��\Q��̉��Ϝ�2o8�Y����E(Q�X}M�p-�b�����ؑt�Ot�<`�,��������fW?Iy�#�Ĕ�w�6*/��xT�!�Oo������P�j�˛�w3�!�g������n�ߙr��-Vݱ�7��,��u��Tx����0-1���`l��\y9�O0$���[��	u��"{�d H*����Vr����3�q�a��)�[�O��_14�>n��%c�D��%*��Z���Ԗ��0a�a�BF:0���]����E9�8���y���'��a��P�d��'��Mƫ��=:��(���m�55�`�ږl0[�͎%�
b�0��y��Sv���@��D;6�f�g�n+��Q�η�X:�1�����k����v ��!![�G���]0 e������N����B�4�Bv<z���DH�LR���u�g�B�����_���3�<���=v���uJ0�"|'5�%�6��ZȦ|]3�����%\Z/��F�eg����>�q��D�à3����S��ۢ^PK&�'����Vח���t�'I���'r���j�zk#��Л �������s�X�<?� �c?ƣ$��m�b�;	��e4���ۼ�a���k��[��=r�D��4�/�WL �.� ������` �Ѩ��䟭}�W���)�"N�Er�,p��d2y%�Z��r�n���d��(�3�O��;��:��!|�A��k��Q͎�-7Gd�u��g�!���;M�+x�1�~Ƃَ���r=xBq���_E��Zd���x`�Jؠ�������eᎩ�si:�A�u�=�����t�Ӑd��=-Z��}�q�'��m_	�8QO
�gbG$�ӾG�P��(�	^"�����v��,�r3u_�ǿ?������I~��=P�2�
~[+9�b瞞�`�<"}�So���>�T�>�#���L=�Y;��/T"����cN�W0��A���!`�v���nJb��v|9�;�J���3�..r�Z�ր8���uÈh8|:F�[��(zj��|�'��#�설B���B�N�7�.�8.�V�@lo��b�T��H���i?ğ>�ހ���}zm�Y2B�oC�&�Tr��3
��Ժ:�艃��G@�b��A�c}�܇N��d����@��(��f��ŶՔ�#9������[���An�&��Ծּ�f�w�A!|�����z�0˛F6��R���e���v�1e7��q��Ϋ�P�O����>l�$�^���ӵI��>{���g��W�)~*Ѭ 6�m�
�퓋� L<C�	ؓ�o���<eC�><=�r��yC�Q&r����߹Z�h���n�ޘВ�3�
�f�
�L�kf��/��4$�-	i�?�d�n��?������zXA���B�l��[v����x���'IĖ'k"И�y��|y���(��٨SE�����q����K�!���P�
͞���[��2G�s�,}�*��)�&!p$Șd�j�;����lI�4L��{�7���lѵ�8�蚛�}�|PŘ�{��&�>��۲�����
�#R^����0t��N�w��:��.3o�ՠ��`�� sP��d��6�d���5$�'/
�+Iy���+��Q��9 J���b_���o8a7�t�ȇy9_�,%�.��	2&��R �WDfxȬ��ɓ7OK��1I�-db@n]y�7��B��p�<tz�"�E.���1�^��]�k�t����Յ虎gY G�tnJ�o��"������i�� `e˹l���da�\,[��+��t�t.��(�7����(2����>͆�����Q�C�<�a��е(�e����K���-ےxǠ���45��PA�ץi�o�� �����|�ĠR]X�&e06��{Vo }���#�-�t�	J?�*��&W������TI�����w���=`�(���Hs�e�5����=�O���e��&P�py�	[k��G�M�V�L῭���e~�GA���?�ªk���u������s6K8�r�R� �q��]� zJ����yK��[��<r�4�h�t�9�N�3��T�&�Rr�+��PO������ ^��5/�r����6t�`��U��Y�#�`�Z���Z�����l�2*�l
�=�)P?��8M[���)P�da�����x?O��O �������Kx?�c���V¹oa�@]���Qo��g�婋��N��S\�~c|AL�����|��5r�f�A/"�|I>-<E�z^Fj��.|�ˉ3�-7���O��=���O7&��������lA��¡Y����?
H���n�./���[C\O�FX <��Y�z녭��T�wå��.S�Rr����4x�E��Ԗ��W�]�6kf<iƿ|W����ᢅ�?�߆l�M�0{��Tޅ�Dh��~%��h�k��Y*��PB�"���I5i
Ɏ7�_qS|6]/<��g�h��oڧ��28��������N�����#�Ջ��Y�&A4fx�a���>*�"�(M�^"�.}r�jb��7�)�Ky�d�0�bz���p��j������p^��MH7K�^�J?�B�9�BJ�D�E ��X��\kk�π�d��z�$��!�g4t[^]j��a�|R�����t_/J'������b��ӕW��ҧ~4��{�>�Z�dѝf~t�3F�I�6Ki����|@ ���z�����9�N���jO�����Olw�

�t�Iֳ*�G�X)��gDq��K�<�,3T7�[pe�0�}��+)En���C(��ND1�l�!s�2՝�.�e2�R���:+㣨�!����d��U>HW�@���1�z�KYӾ��=����V5��1M*�1��s�y��ֵ޷���۝ipz=���!;MC�,��_��+}hul��c���̻5K�����[���l�`�Qs���7g�hy�8�O��-l���~@�y�=4�k|��f���}���F!?`�+��h߁�Z%:;r����d�DY��v�q���������&�ǻ��<BI��IBc��B L>�U�>_�sbs�̊	(ϻ��j_�/7;d�l�����U$�
�܊s�Ƽ���aڝ�-�a��!�P��R����z֊X^�}Ⲗ���W����:1��a�K�9(�	<�^��~�5fR���E>�F�`jHlK}�����0i3�/NIx�&�-#��
,�:��\F��?�\�~�xl��2&��ݳ��O�Ig�a� B�p߇J��g�_	@���d��V'Fa �n$����"瞚���s��F}3տ���ĖKV�d����� �
Z�E�m�(hN�^(:�X�����k�(���i��2�X(Lc�9�A�@*�57���_�(�3�3׃�X�;TK����=oU�C�C9��'_J�����b
1gC _��脙O����9� �i������dSP�9緜?��Q�0����!���B���}�n���q�9�R�m%f��Ӆ�΢~�M�-j�a�Ѯ%�7�c'L�a�#����U�2dih�X�������f]���E��oxf��1�Yg���Y��o+'���_�@����eq�P&���1^��t���,�"~�'y�@���/'[c�UL�L���U�7B(׸$= ��x��݊;P����`�?�[X���]�'��}jV|�M���}����e�Z��}$�=GP�w���L�����t&֡}���L���{}��l�c�r�xi��gf��nH"w�qɝ��|S���s<&o'ڪ�Jj��S;��nÇQLyM�*k�""0�$HR��r�1O��lOՂ�-�2^��:�E�St�=��;���%Doo����{���k�^������l����;�
���*ʜ�������>�gDF���j9f�oT��,��7s��9�@��~�;�ef�(�	���j�F��X��|�dҨn!�@���%���դ�����E�K�� 4X
.��d-�k# �S,va�E����6� ��iVZ�	,�	}z˝��������x[qB�I_ɶ��}I+9'�9y?������О*���+:q��X��"�l�@�J.� �v~ �Q�}��:nǹ�_��j4y7��\4��o�7���9* Y�$LyGuG`�M��򚆗��iYp�yUc���lJ6Cx�(z���}._bkz皮���ɏLG�=�p#�_��Y����r����Vl|1$O2�I>F���5�b����OK������R���-M��;���4}ӕ������-��5����?��u+�}ezB�zU�"����5AK\�\L�ઃ���įlWh��u��Έ�<�U�k�w������8Z7��J�.�2�;��]���;��<��e�ʹ��D�<� YPw�`��o��z�`r��|+C��N�R^|�͸���t�P�Z×o+�$Us�G�{��f�s�����7t&�ѤkĳC�dOT A\Y��lMlA���*ڬ!��[*i�q�v�;p�Çz�W�3A�9/5Ch5\C��ً�ժ�AWn���^9����\����l�5}oxT2칶jOa��-�",S��?��n��3s��~�K��z��@��Y/��^��z,s0&���}%�}I��W3��t�l��d�h-�����l8j�`�TL����Cb\����u4r� g�ު����/ G?��m��ŗ*>Z�p�9�>/�ޠG6�9ǡ�"�F�1����/"��cp<�{b�E�}G��0\V�X�=��'+dZ�h��.<�z��N��g����h\��G>�lM���F��*��:�S�W��#n��As��	צ�N�Ĕ!G(�9O���N'���B����y�Qy���|�'�7���П��Y��~Wt-F�\�����x��s��ނ X��B��I߱�i΍[o���W,��/J����廖d��s�ĺkf��)9P*����r���%Bȩ����"�1�L4��?e��$s�|`s`O�L�WΫ_+���鋍3���$'9�KI]�$?7�(�t�S��-��EBc6qnyZ�e��9�.wv�ϛ�h�p;�Dv��l�Ls�Gx?����Ċ�j�'#�I��nw��l���=_�x�gn�~C#CC���1� �d�R��>S�^��4z F�i�Y`G�R�y6���βyXY��n.P?/�d�f�u�Ċ�59
!V^WTT\�)������%'҉;��bxs@���Wֶ:j���Ї�.��
RKTkz�>�G����Ƴ=��8a������&�'�Bgo��2;�R�*Q�k�wU�9�bj��h�o�T���~�H�6{��H}Yy���^n����.i�T��/7O[8���;O Y_	d˥|<�f ��w6,a撹�J�q�@��9��P6�4[*ER�q` ����IyQ���
��Ԃ.�3��<\q�e����^�1��xBP�d���s?zP���-S��D؍������<�x�iqJ�(������Ym���l|ߪ?5鿧u���L��KT�IS-��?ƍ�BqU�F�x=x{�ã���t؝,�|FlNz屔?�'$�U['dcy�R���N-i0�\�����j�PE���T�b4�X�@ٙ�
,v�;<�j(�g���?�qQ�z��;B"x�\"���*��߰)-h��V*�çXڬ9�l��Xn���~|�f����iN��3�\��7�b��h16}�s.�у�s�z�֕�e2Ag{aǟj 䎅�#7�U���s9�F���Cq�"��ǚ�l�<�̠�d�b�W@�e��g|�-p�!m0��jMC���0?��Y�AW��������I	���Y"�t�FҦ�e�������9���.\��:�
|�+ t�M�ɦ��E�̼T���Zd֒�j�`�ӷ��Z�m?�������ZF&�M��HގZ��!�P�g��5-�bw_�*��٤���O*\�S�J�.�D���qQ,�Ċk��(��\����G��ګ_q[;����U�P��iBO���\���D�Yo�;�t���~Q�5�Am�S�����J=j-��:�Lq�(L@�5u��L�p�Qܘ)�=�����	��Rh_#A�7T�ò_�~�|�gUڼ%K�o}딬`~�z��>�(�#g&��Y��@�T��9ڎw��5�l���2����Y�ө����z�#
ßs=�x^-ᤲ���B��W��F*9�µ��_k�{I�@�gd��Sx䏀��WM�
-�5aw?w���|Tآ$D���ǧ�5��~�����'��@;
���W�0�q'qKP̳��[m��(���өT��FN)s���C\{4��Pe��$P�������b��H[�WE���
s�UP�������9Ǧ��cū��&k�a� a��˗����%�	ưm���|J_�J�-L5�SQj���+���AQ�m�i(�qCU$���V�et���hy�����ń�#����ac�������</��I��7���S~I4Fm�E�U�r��UDHWr/5Xդ,iu5�AOL_�R��q�nD�����Kr�����C�[�E�}��C�� #����-��2(�))���A�F���i)閖~�|�Ϗ�������^k��u���9�W3=b��@S~�6r+�B�����$?J�.��;U6^a�jǽ� �����¹��ZZZ,c�f�	o*.�c�_�G���ºɔ�>�$E��ajG�֯�z-I�:�0G�ȈLV����)٢>�<a�%��T�Pg����ఠ��qܪ��m��c��xPN��\���:�h�����]ԲiEw��"q�������0����!Xat��j�G%�T,��~K�=&�~�F���%�5J�'�h�J�fHw�ۡ��~� ��L%��$G�?�fk���$䁱���{@�f�.���ǅ�O��FF�����3X��Y�TTx�>z��G���}_dÞ��)ۼ�����Xh`X��o�JT�gj�������"xܽ�]���9᧡���o.��n�|��{��R2���}�R�������-,�0�5�٠��_o�0/�T�t�)�¹��H���Ĕ�r
r��4�R�K���h!�~����@d4�wvv�G��&�޸�t`©���$5��bU��j��Y̶�(;������׹�=W���U���m("�6�t�ѵ�4I�.�;E�\HgN��m?��*�� d���q�[�W]����B����D�"b6f*p��Bc0�ƮL'l?W��6���DB-W+�Qn.=���r�D�G�rq��QVWd!�b��8ͼ��|8�!�۷�����x\6�Y,�+����w�`ܔH���YkVjrr�A�f����17|�+�gҢ*,��SR~��!Y�a��y7<�����?��l~��2��U1y�M���H�3�c��f�g�D���i��`��Z�lTQa����o�;�T�V�D~.��S�%��iog{[�#��A̔ �{
"��e���In��i����kt���1��/�2ĊJJn����]	`���C)�oNw�h^ki�bx�f���ҹ��*ϘXo1�We5o�s��s�B���2n��lRҠ���+��լ�͛dE%�k����Y�X~*#d�KJ�ܻ�!~-�RRRi����<LQǱl���gKyT7V|�7�a������MsS&S�М�܍�A?0�Ē�QW���5�k&�u����3$$$���
���(3�}�'�Y���S�Ǵ;$p���
y��߲1���WU%�q�����_]_������'ZJm(����񋘣�`P��9[B�~���M#
�f��Z��<f�֋E���GN$���S���8��2��PG�)-ݳX �+��dT��{���8�Xk!]Y�vI���/��[,�D�e#HB���z�͉`M�$�ð�H=ruEIp\#ll�8�f�Ғ���R(L��#^�K	����;��O1_��)3@������*#�Vj�pG�@׵�h�^�芓�3�*�L�+)y�դ����cD����D�Z�b�ϫ7c�,QO��Y瓰��b��c�xUx��mt��O6��˯U�{������`H���<?=?G0>T��tl��1H�A���B�w��.@��}�����N������fL9��F��������AEtIIT��4�4:�Z�vx��@������f�C�2V7$����W����2��Cڗ�����^D=��b���+��� ���D_4�Ћ>1���"�C3�i��+��o_�ǟ���ӭ+zMR����=��K	�f���m������������/_�\vJZT焇~���������H���^A1�ܾU��x�'���kɺw<6�sY�jڥ�L�lzEp��Fs�0�%?rDn�"�6|����$V��Gf�����i�3��"�s䙘%��A���?yn.�V�:J$C�Ss������Ї�G;U~�v"66V��ּE;D��b�#H�d��{*	_Ja�o:�\��Wswf�P�nn�����<S�jV�����5g���׬��Z�u��	B��O� ���0?p�
�1xyy�EM����IO��DQF�ujKh�b.�^��K�4���ᮡ����T�}Et@���v�n��y��|���Ъ��2���F���oѣy�mɞ<ל�9��e!��ΐ`hh8��@��Ǳ��t	,i�5��:������w�o( �q�4��=�l����G~:�E<A[��SfM��mo���c�2]�<iH*�0d�r,(��&��AJ͟������#jmc#x�2�b�O�FZ�5���ϨGF@y��ʱG��pA޲�X���M�$fR����&{����sn�8�f�IpS����N�43'�;e2211m;oCȻW��σKJ�89���҉��IJ��2	(}0���ι*��x�b���g��G�ɚ���@�U��9��q�T�Vt�V��J��e^�uE6g��D��������y�=I�t1gPHԜZ�f�M����N�x�cY���sȼ�WdD!q�v~�e�"g=0�����O�~_{c���Dq[�����1j��5}O��n�Ն�"�e|�X�Ʉ���I���L��j�.�:��J��%V�`A@�N#%fT8Y��:Њt8'� 9iA��[��3,���TP*�R�/2\�e�)�8�%�n�(L��M�[O/���J���&����H�ÒQ��}���ϟ�ݱ�F
�q*�͗�󙉅3�;^~?k��\$��;�3z�]�A]Y���J#$�V�<��`�ZF����G�m�`n*-�.��͔��6?=�M�Ud���h��.xQ`�$�Љ�z��d����"� C���_�=>�kt��K�E4"vzz*�Ljj	�_}@�����f�*��TS�H���b��U�p6���P~
?i����� �s7&{���yqZ^^���E��/���-��m��@sJ$�i��`D���৓v��&��]�?����HI���s**����\(Lf��c���ܞ�� Y�aw���8��qw�G�Ak��B������_J�GG�j���n�G�5HQ/�Ω��a��'�-]��%��H�50�[�[��.6��r`��0"ĳm1y�\�.߇M�1\w����D��v����tQyv󢉌����ZE�|�h��}��G5hH�M�,K[��P�]b�-R�E���ڰ��v�3�^�Єܶ)����x�Ù�]����ȞF��O)��?8p m�h�F�e��{�P�Y��j�|�(��EK`�	��蠄N�]r�P�;d�e���OY`�VӟQ�����O����\��4m�L5Q��C�/?���u�e-N�˓�:l�X'3y��}����E��b)�����}�%.L�t�m�Zq���_��Q�|_��>t�*�@���O�e����)��5��O �Ȇ)���[7(��'�'��6o�>�rB-޿��I�R9c5��D�4�V��6~V�|$��$[�9r�
M��d{w7@�,R��)����z�!2���\�$M&ز��"�I�A���W�P����)-.�	��x5w��i;˾�\R"����[�����jsy����JPMI	��2�x��ѵ���H�+��g�[\�|��N�s�� �_J�А�ʛ�SB�0"�ƿ�%ł2��F�l�����>��w�F�g�%�1m��gO`��a��O?bS���8}�)�b�����+����Y��
���3?ŘQ}�Z�]/z�f~H!��;azc�%t��o�8��X�F���R�y_"�c���7CLq�Z���NRv��""����tp|3)z�D�iMo:7�GWl?�y�BgJ�����|��ͱ�9��
����c��D�a�b�?�������n0�=g3�y����%:R�eo�
�^���n�K�	/�ȉg�t4��$�n�m$05J�����m	bcx�w�H�T��?�V ��BKd�,U����t����k��!�v�(��`�1��]mc��Ӥ��~�l����Uhk0%is�}��
��l��i��Ą������f��weUՑ*��X@�@���[Z3|���W����Hd��/`�ߝ3l)Cs��b��eX��㸕���\Rr����a�OVNn�L��%U����S΀Ĕ�kjjZ~�D��՟�b)N8�и�Yj,��u��̊�D�w�Kdt~�W�W�3�̠�jVa*�Ԯ��NT�h��҅i�W�ag5߾�|oBN�Ѫ�R��W�i����W�Hs~��G��o'�M[���禩��*9�Ƃj����	��̈́<������K�[��
`U��?6O$K
[0._\綴P.|,��7ŧB7s��t1Ml}�*ݚ��g7{S|��$��V��)���mf>��N��"��O�~[�����GY��)`W�褬�;���z��-O�@t�I����.�������Ց��4언��@*��e
���R���V��l�D��NP����
���Eb����-�x/��jO0S�d����˸��ș���-�_"#$�Cπ�E����Sŭ�W��
�\5B�Y)bw(y,6r�����k��fnL�@�Ј�47�=Q���~Mڵ��jt�o��EP9���%��#��߽���Ѷ-�$�Ÿ�	�f5�(��8Ŋ%���j_ϧU�>{��I��*�
�5�l(�X=6#��%�0+Pj]pؔ�`��wXS�u��7��U/8x����Ii���K��U��M|� ���i�����~?Zv:h0~ӫ��l�@���C�n�5��ޚ?���U��f3��rvмH���Q����`�#��� �cQK}��'
�.}�y%$&Z�������Vy�w��k&TJ�UI�� �Ѩ�� U+� ����
�!ۡT�}}h 0����q��{7�����޷i)��$2�c)WWW�<̈́��T=v�[�����#�G��RTIe>�>)���CBz���mD_<�q��O<99)��|7h�G��}V�����;����� 27����v^0Ȏ�S��0U��Ib������ĝ��UA���6P,�T�VCO'A*���y�ЄxQ�x��d,t���))��:[�?�'c�2�:U�?5�MIA�_��%��2�Q�h,_�ߋ�-�����L�{�f�{E7*!r��̑u��v���O0X����νʾÇsM.�O�6_SDzf1����IH��7|��|�
�Ft�R�UA����K������qW��I-�aH�U0�G�{�m���wo�d׹���Ԯ�9��\�ǲ��(����`A.�YǱ�C��&�{����rq�^�ɚ3uo�O�Ϊ^�7���TS�{��*���#���ػS���TX~�=�ġs�9r���TMW���ٙ��Z�ڜ�F��+���������;O�7�9�%��	��qZ��q��8^����"����>�����X>�	�Z]R{M�Z��2�M.�h�].j�s��2W�:3f���t4��ڊ*�(�Jլ]ݴQ�_�X� ��RH�����b�/��G�0(�r��r�Ѳi.���Q��^��
>%A�B`?�,k!'����y'�����A;;;n��&X)EJ��w�\�b�e���P'# "ڭ�qi���cj�~�Z��a'���p]as�,{�E'%�H9��d��X�T��?`�Y~@�{tx�Ʋ.gVu���|������wE��C�Sl�C��FB93.^ �[��O=hu�t�ȳOcu9�U�G��Kfqh}~���z��
�o�aaa6m�?����C�1�q��$���wd��UT�XN]G�q����//��o�@�^t�I�lF�+n�(f>�3qݦ�z�74d���f�LRF���	v�/>c�o�0/	-��!!nd��ǃd|I����󑥀��3i�:srJU��iʒ8�)Q6ś�?��XY�5V$�e}�
h�#��*�8>��[���%L�u�5He6�W���~�KXXXhd�X��;JYY�=}�s�kd�A�y�أ�������i�wn��gI�1�:)
��4�m�0�?Ez�R������Ɯp�ǲ��E�h�#+���J\8�<q�����:3��y;_3YrS�Z��C�:��P��}�&���^Л���l�8͒�0
��t~�4��!�2�u�&�樵nJ�м�'�J��5.���^������Z��������������p�e�X,��
J�����:8���'#�`k*Rlsm�"A|�c����-�Vz�8��#Z��x�����}O��Ϟ������/���Z<=������'��U7�\�����֚/7�.//�)�zOD�V�)s

~|>.��GF&�����ԕZ;�������=9t9I��z���*�~����5/nHHO�������]G�0PsII�]Gss3�."r�uك���E�ժ��`B�[���`yצ�U��\�vQ�b�ذ�J!+L~�D�<>~g%%Rju(:8hY�a} Uءe�>#*
׹���p*�Ŷ�}��c�m'K�P�r�:S{�	���~�w����;����q^e-;��"	̜�<=����l�d~ۋ�4*�<����±�+@X?�☿p՘г˸���ݭ�)b���z>K�G�^�g�knk��8;:����+ P�v�����U�,�u�X,-��������N�"n�(�r��I^���iW����|��5)�x�>�%2G١^n�T)�7)c�}������\��}���Sd
�λ���Fl���v*�I�������o��ڨ54h!	8J'e��_���f�IA*/f�U�,����N�Y����c%us�h _QP�ˋ��W�s��-����å�Db�|�r/>��l�E9Cԇl�s���Oԋ���<�Qy� �_n�[��n������t�K�����[]=��i�C���F��� ����y��iii�1�]Q�9L6?����OL'����y��f�o��"�K�վD��̭�(�b����˼�/�U�%Z�	,R��"�b\���ʼ�TF������ ������=��X�!��М�C��ҕ��e����?\@M���</�Ɉd�a�����ѱ�ktZ1��A���ɨ�����+Wż��=K@�d࣯P'���Z+J����ֿaL<�!t2��r��)��ȟ�ru7�;���*�C.W��2����H���O*��P7g���އ�X�<kk������}Q�ʽ��(�Y�#$r]��8���JW'��n�,��\�Ʋ�a��1ChG�T�f�,K�\h�ϟ?W���߂U/��)���{��`��	���I�w�{���h����D��8��=�z�:-M=OC]����+pe4��>������dnnf捍+54V&��݂�tU��GQ�ӡË���̀�~F� 1_!��_���A49ǔ��!�{̐��БM�~�y,�!9��d��H�0���Dݹ�w׿����7g]�����i�����p��nllH"�	Cf�=���iE���H�H0'�R�ƾ��Oy�b����Ƭ�X^�L+M��;IIu=��e
�/��E�?,v�W�tb˦yLg�2JR9�"=z���3���Yg0V��bU��C"��(�id�k��pQJew#%'�ۦ����k9F��}Ş�7gb��<R�p���߭���b�~���x�ͧΚ���2�����
����ʾ�}ο���T�,�z��O��d���7��y��`z�!V^Qad��U���y��ߞb������Y�((�o���ų'���H�j��[[���ަ���x��jͭ����G� �[���ot�e7��/=�w�y
�w����5�[+Ds�za�S0!�-!������oooŇ��~*���b�k6�4�f��G�/80WT叉>rr$�(R��taa�l��*yZ�t�P��� ���$ث"���|>5�pn�:cm��1���_JJڟ��p�>�g�i����|�j�����H4���ݰ˓�yˡ���v��ӉO��#'{Ijbcl"z6��<�"Pw��!�j:.�㇡0���|��Gq�M{���&W���7˯*C��ͮ.�Ac����f�@:h�
|\2^�Uq[O�D&yߞn���i�+{rN�����%�� -$RRR����B���c�ʊ	��Knmm2P`�T��Lb��KJJ������+�}�vk����<@��L�Ϲ]SN��������H���/_X��믺�el۝��os3G��6�7S5��Ҳ4222m�0Z��O���k���8�G�P��͠�KO'�˖��8�XM��'Y��:4$hR�s%�Q��h(L��:��Nƕ��Y{at��ʳ� ���vo߆ ��>^���D��eC�>�	��;/�&*�$&5YBj!RLt��p�8:����w`N?���߲��P����������|����ͽ�h��%č��9�)|1���O�J�F�NW�B�O�[{>q�4��Qſ��hq�|��U�
�?�����oMϘ�,%X,�zD�FG+n����,�:�����[;8��5!�ș+"*q*��=nm}}��h3|s22�7t�o*;�Q�֗�榩_B�>��
��'���f�܅�X�B�i�Ĉ��3Lhn��		�\[��iz������5�V�(�r�FБ��֮�u����yi��$�9����"� K[����gm�?���p��xv�x�����4@�J`�)8�ssx���w��ȇ̩/��~ͥ�A1���b�d���W��-�/ ���e?}(�/3l�����SQ����).f*�gcg�B;pz��.X n�)����yYY�
�踫��Ơ�@��
^(&]h��<c�gr�e�!~j���PSC�s$KTox`�d5�w)p�ɐg�xq�D��������*��\1��q&8�����Y�9��f�����/&�ʅj�J�xӉ������|�枹M�]�.�D��%_���5�����?cW��߂q|[R���MgSz�@ō��X|����tP��Ui}=��B����2�5v�G��@'֕��;�?Gh{F�H�������[��$R���q2� E5(AϿ��z�<��" �o	#V��Y��G'�����mlm��.tӇ,��K��[�V���>	��:��g@��ƥ��\2�ZK���5_���,�?��^k��*ϓ�!��<�����5j+×Y�0��Σ՞ܢ�p6�Fؠ��EL����T����Dm\\�hK����3��G���JKc�AH�����f=��5%�l���pS�T�?e>�_O�9�lM;�?ҿ�v�`�ֽ������cOH&��S� ��mn�@�7ekr1��pe��L�� 7���M4	K^�Z��>��o~��Z�S�c?�x��®[0^>�����ՠ�9ݏ<Vq�)Zgff���������4����å����D@���i��>��%�l��a?;�Pm}=��+��wɎ�I�Ch쭋����1.[����{�D���Ԟ�>��/s���3K�������?��1=u��2�s�󻍕�.ݾ�>��]�������qq��|%����O���fp&R

�,��}˂q����{�5c<V�̛Ùfc֮��[W�v.�h�(N�����,,�$L�5������|���M�x]n�Xo?��I>J�5������-��҇�=���~��VX�H�O�lq�o�4,�?k���8@����l���(�cqt�g5�<X�pm�������g_�(V�hnbfe�:yL�������ir�̣���}����,��YLI��-��H0r���.���S.q����cY�� v�-= _]<p������B�z ���R@�ڸxl:F�!����醀�Z�R!���0���-���F(�U�rO8S%>X]�8��V� � mG`A�0հ��Y�'��/��������;շ������d�M���%{}u����a5�0������4��2F`.���N�[�JJux:�0�X�n@>�M�|��.hX�N=h�X��-�d"!�����6ud��3*��BS�v�sa�+'@U�P��5y�S�&�ZJI�������%�������n�����v܍j�eR��
	����ab``4�\�n����.[$��$	5���h_� ��t>[55����\HB��O��C�Y���$�b������b�6p!)Dk��ЍOs�����{߲#os�rڂ90^4.�T�^m�Ê$��R�J�7L�w�l�d�Lו��tY�n]�&�jqQ-+�~�ZG&����՚��Q�V^_J����!�pq�qH�{DF�j������I}*ҭz7��t₂P�����8��:�b�h�p�j��Hкޡ!���DF����,(}i[5�?�݆͑��E*�) ����vQ�Έy��hI]5k���/S�sJc��[�xJ�U�/�A~��,s��-L�i�;�F�ݩ������K6`��P�M�n6F�E<+���QC �A���Qi6�y���6 �����F~��I^���NI8 �K
**L�u��!^7�"�bu�I���	睋K���X���1�n-���j$kN����3ZV��_�n�V�y�����|�8Y#a�>~��@`��}�RS�b�?Z�(�����:Bo}��O�p&r~�Ohu���V��G�XZHj���immm[W6��ݽ<<<|����\ټ����'K���G���U��T����^ƞ(pg�L�L0ݫC6�B:(:H����K�j蔸a���у:z��$P�0C$�)�cra�c��"t�2����E`�Oٸp��ut�lq������V?��z��I晇�����Ò/_��x�g�ށ�s4�����$5H�Y�e�4mYZI�6szCDv+k�]�:��(��J�׍����ec���\���xK�nrխ����
]��tB���Zs@]-
(.`�7��� �J4ōZ��q����t�zhD���K@��3r��3��!���k>���I�th��w�T�[q
\p��|����N��f����(쭍MЈص�E���A4�M��d��Y��A��gs�-��߿}�FN��O.�,�0��$홌G�Qw���-h!'�|l.��)cʱ,�7�|����*�5�n�M�8@�⨅�UTTP�^;;siik#���zv�̔�m:� �i���lM��Ke�cI	쾥ȦÙ�8����c(l�+K>��5�9J:�����&��V8A��⭭�� =�4K��We ͘��e�~~
H��E��>~�hY��h�qy���Ш1�<9���oi�7������dWϧ��ݵ�^��t\�M��w��PN�5�{* h�����.�OfVkϟo�g%�F̮tE�l��s���^���$X���٧<8�=�D�s6�م�-��� 9��\_`�Ǵ ��1�w��M�F�� ��fәH�oǢ�إ�v�?�+to}Ƈ& G�U��4D�
2��;�������~���H+*Qoҹ�����̲N*HNU��� G�o��8��C+.$).�wu�:`���x�<��Kf1}�W���璒ps�;]7�3G�\i�����ce%��+�n�{{6V���@�`����x;ɚ('|~�J��j����@ )��Á�*(���؀�a�a��#v�sA Wg�����~\��7���r8�׷ұ��{&8�m���g�C�YF̌P�%E
Z��^,��!a����z�MO�$������͓Ό�.ƀ���U\쪰DoO��ǘ��o����[Z@Z���A�2}|����i��)�k�|{���������쑓V+g�-�(�T�K�4�u/��j��,�f�P�u��/Q�Ќ�=eM����������8�s��� ����lf2*E�ݎʫ|U��ٗĴ2���������c�Cr���J��������R�"�D��"������N9����67� R��r�%�-{Sg;8vFǫ1_o���dH@���ݩ������_����0i��69yy�#Yլŷ�$T�{5���D�z��	-F��>x�(.nԴ���v��h�ԕړc\��5�fLkO��~bK�����\�TIY��cH$�B��k�!qTV'�9,4/@�z@��������h�y�����˂�l�!�(B��}���BJN^��<Hς�/1rDa�Ҳ2��ˠ���Cf��.���v+����rf�cb�⏏���C����G�Χ�7!��,���`�7�AS��b���*�k8��ia��mw��(�FσR��ot�ѱ14��U#�_�����k"�5a�����!��X@DHX`UJO������il�M4�@m+�w�Ci|�`���>��������������Ņ���:~nd���H����F��<����!��ӗJ@��ht�CfQyo6|�<����� ��]��t�8I((<x��1�%|�Ͷ��|�l� K'��H�t��I(�-�	,�^uS68�n<��-����љŁ(����<�;A�����,���l���63[�FI��<� mE�Yp�����D�.u�[�uqz�1�	 �a �k��U��Q���;��]�^��rsy���;�����ㅑ di�M8iә�����:��DO���J���vMNM�1@nL��n�Y��@�i*煹s}����ڲ�C��o-�����-�1�_��b�~[��Bl�Ě�KG����aJ3l�������E��АH����5/.(���I�͑����>ќ!$\�f����-c[��3Nd����]�s�)��-Sv����Im嬆�"ܕ�;*}m��0���	(���zAAA�����M'}Z����=O�<["FVkc!)����O���۱{�3ј@P����������q�����v�zܙ�<��Ɂ >Z3
��0�q{S,{$����b��I	6�!��4H����s����C���o����fk��}�u^lE��!ہ���-RI�8�|rٱz����G>_[�u��	bO���u�(8�@\�%ft�^�00���:8���_��{�ü��cx~�%�|u����
N�	�9�&$"Zz	z�R��3�Gh��1e;fĘh(V�<����x�4�{�(�u��� �C0�ѥ%���6�G%������rr$1D=�_f��2�Pŀ��uzn�9����ȴ`��CI's:F���-��L��$r,�ET}D����xAT�s�4��]���ђh�k��y��GIt�K��L�{�E����㯧��&������-��gR�Խ:p8ꖝ�����寧��Ԝ�+�Z.!tH`JJ���5�⚩}w5!*���]]{v�.N��~_bիߛ�>$��2iY���~N��X)���Q�h�t��̽!������ӽ�C���[��q�ys�S�>�	Rg�=���Nl&:e�봫�2_�j�����P4j?U%%%^�����,��y&߱��@�H$�BƩ��@)�W�����?5�=�\��A�����[���SW�SiK��/4��P�;��Y;��c�o���� ���yP��wG޲wbd�,�K���JJ��lrJ�3G����B��2�ʋ��xz�$�<~���6��Z��vv����l:�����5c	9��+5�5�6C�YiKߑ�@���_��z��O=U��g.T[��F�g����#��7K��r2�(o=9N=JB��Eo��X��P9�m6����w�����S�����ë�]#�f2^/����|á�����1��j�_͖���k*/����,��B�?���V�y}�:��A��7ߍ�OFl:ա�^��O�{�c�V��w�+�������l��R�IW�HelW^���!���CP`�O��?�OGo���͗���Ѩ_ˈ�n����u������=�zL��8�8�7ͮ_�K
ec-S�t���[9K�TJȫ�={i����gf�I�k�z���6@�E�Bi�m>�8�C}}_�����D8�G̍�fJ�0����wvv�'��#M��X��Ie7����d��y+�F�hP��2K5��:�t�l-��AYKC�˳�@���k���p��4j;� �&}�U�H�'	h�h\IB�|�!U�kn�u��e�U���
�Qǝ*�k[XX�{��yQӂ�R��?��Q���~s��ќ���~��l�rή�8�P��%��l��.���o1����������ؼ�Z�4v��Q��� F�7���V$��8��Wk�p3����zp����߿�G��N3a\�)�|w���DF��i�����TW����P��;� 4�¨F����,��'�[�����G[���V�Uy�f\��`TQ^.f)����4�� ��?��݄E�~e)��:��'�HFh���`�nE��DD��l�Q�r-)�8�:Μ��y�f��[�6/}�SƢ��& H!��d�Pz֩X����_���@��)���'6��۳�N+��F�a�VZJ�������՗t�{�h�Z=c���Wcʗ*M0؛҂8s�S��ODt�̥�u�+�Р�<�S�4�q�O�������%�1�U������-��y�k~a����˞�ⵓ��DD��k����"����mWE�-������@=Y �����LE�3�Lү�� C6@��5�:^{�tw��n�*
͍��	3;\l�����&�Y$���D��Q̘�ؑ��󋧖�BF��g��<�6�����T�X�S�*ՙ�qe�<V�����" ��ip\r[q������I�;�7,��W<�l1�{���4�������T�%@���s@���r���{\�:Ć�y`�{�1�5�}���u$�k\�^W87���fL����!�8��٤���6t�9;u$m�<o��߭���)3s���Kh.K�Px�/8f���V�n��g�T���NLo����S� ��u�w���b�cu9������ͬ�����yy���E^O�zh!��*�#P�u����������Db�K�cӁ�%V�� `�5�	{K�����`-�>z�ش�2ϙaEn')�Wm�� ҈Y���=��e\�I�7C73DR�e?C�cx�!4�輺�����j����f���Ɵ�:aH�qbȯ���V�[JW�Q3��l����B��"�
a]T�^S`C�����V�z�G볋x�z�󴨨�Q���aB�p�n�=gv&��[�f��Ў���[kkk�� Ҏ	���׶}����fGe�x�&n�:xP�d�������ͬ�]0�lV�f��qM;�&�����F��?�<۝9��+����ē����c�LI��3v���2AƜP�RF'&�@x�f�U�==_�?���z�F��~�ZO���X���R�}(3	��]� >Hp�)�PL��o�g(}^�:}�I�$�C�A�>rrr�*��̷z�@��#�����@n�#�3T�Q��^7�;C]�u�{\���` ��!h_
 2�˥)ۍ�R�{j>���B���z��x�~����
���L�����TC[A��_����]&�|��ҊW����i���-}z`&[�S����e����r������5�6�p�s�c��V�A:8 ��åÂd��� lH�z¸.�8������p*�P��c|�������r�u�A��|'�J6C����� Z˂*�9�Ө������Ģ���^��B�͜m�k�&uh��Sw;I��*�$�3 l z���Jp�y�j���r�/~��,L-.�q�l����pTb-��ۇu��[�~�u�@�98.���,��	�|"�*�04�����+��� �%�XY��dv��5'������C�"�P�b'����,T�l��v��\���q��4`j_��%S��$:�$2V�6	�;	:�1_���l�'�x ��s�CM�u��7,�?���h���Fc�_�PZ�d>���sh��sls���11}*�9��ߟh#q��#�QqT���a�|`��Q�=�X�����F��N���E
H���)D��䔔z�+�� �������ʊ��ׇ2�������(�)���,�үa4��*ZX�玉S�mA�͟��.�M��]B%`}�k��B�,_�
�lE��_h�z.94T68Pק�?��}��-v;z�=A�Po?��\��ƅ C.����&C̨���I�8��U��Ȑ<.�:���vu����t�4H��x~xwp�M#�����ӧ��=!�����!ψvP'ƀ�(7hq�K�5Ru�ܚ!a����{�¨�t� ���a�0���S<Y�,�����P��;)I����8a>�4��m�cɏ]b�DM�h"..�ݰ�m�9�?t�~_m�m�}2^^^��F��?��x�n�&�]`��ȅe����?<��X4���>�L9�8q�8�y���%bS��Qlf��AN�>Kk� ��z������c���C��oo���;Jꉣ�Y�wO%''�c��Z�L 4N�a�z���z�k#������ps�(�b�QQP���D�A�[�{Z�z0Dz�%�h�iO�PN�D!�=�7�Ul!���Lt	�;G��$Y��Y_�� 2�7�^9�CjiբA؟���\GD/j1$~�q�:]`�3dccs�"|�gg��j4�xq��&��_���O�\_�}��B<+b�e��^� �H@��[)J	�!�P;`�Bn�#��<���n�2��[��hh8xuu��G6_QPRޛ�V��F[��J
C���,�|!�wu�K¤Z�l���%t��$�v ��]3p��;_+�+���p�^*�C}�{tc(�͸O�����G$I;`<\\n����Oq@Ș�%aoTT�����y���1i���B ���C?}O�{{�!1{�RjYY�8;+�)�����<������Ca�=Q�%�XT��OLA���
z "]�h�'�<j���:Q��u^2[`�o?.�����<Z���7�*H�S�E��1�x��d��e���w��j8YZcp�2y���C)�x��rAA�>yVs�w��VS�A�����"��y������AM�]�h�B���"EP� �"�H�����	%�J���"���Q���K�Dj%9�����?gμg�3�o!${��^�Z����PQ!���Xt诞7�
ԑ�WR��<W�������(~3��� X�m��� ��dtioR1��0��ˬ�Nb:z��Y�A�E�z>VȢ�BAn��4t'��VF S!�3�Rk=�_�& gIs����!u]>D�~~�/d�9&:�UNN�d��O���D���0�)�~AQ11�fG�m�>���}��wE]e�^X�7��/Sc�d
#n����=�AM�I&��T��̨C���Y�7�}�XI��݇���8�r�ox>Q�����a^��T���-���M\�ຒB��e�B#�ʆ��$=�&�v�2p��O����4���a��3a�S%\� ��������l=wirq�D7cF�~j�'����pZ��p
E �X<�S��9?����u��E"t>z���K��DM�=9����:LV�����~�� n���pӲK
�]�v9�ש��刢b4�i#\I����#쐻�?���#WG �>�꯽{��2h�Ү�/������'��ё*�	`ޗ3C9��v���
&�%�L�x,�k��tC�˗/�_+wsut���a��iR^�ɇo#Y*�7����k�&�z���.+-U��aH�zg-�F'������z��w�����)���S�(
��a�`������S�@V|�g*Ć|{��~I��e��-�xDC�> }%�-Jy`�A|e�������P/Yҽ-̌}��<$ґ(F�FK���OT?9K���l��ʅ�dw���TVV�H;�<�34LL�]:yU���8iюiV9�6�?y���@�N�;���[�&k�s��jIⷤ�hg��[��6fփ��nQ�lL{?+�sO���m�|`�`�>������WTlI-+)�\Y[�Q@�{�RZ|n~�H��&۫�{����Jw0-������	�1����7�����m���O�,�Y[� �'��:�/_i.KR�9�����՗w��&��7K@�:A�?�|�z��'nz[3:::`|�4Anp��i���W����ia��h�{
�c0n��~�`(���Nq�ij��Wl<�
̍'������?<l),�ko	�x�(�
�B� �c`:M�4ed'�������uq�Z��O;	��(@\����Ǫ�7�_��dR���{)a�թ�)�X E�qkk댼u�m@d��ō�՝�7Ww���M���b�J�g?�����6�$&�`ݍ����L�,�;M��ݼ�
:��ýLI�nkB�����9�5S�&&&\��JR]Tq~����}f)B}��H���H]W�8����F�P_�"�HYjj��߿o���qD)\�C�����g�d�x�x���BTDͥ-����.f_@���������"G�:~K��t�@,�Ib�`�A(�'�e}<��0�ddi�P�t�Qp��@���o��/���@o��MC���r���ia�c/��OӯF��}=�pÈ˞e1��]�̟v�1WCC����9�����|F����îx���e`��ѧn�
u�v�~������g�oIJ"̽��,���===�m�a�k�u�?��1t��G -�^ziH����w0��ggg���]��_zP5	���X� ���������w�|���U}�H�*�U�zX��gc��ڔ�]~jj�����FԈ������q��UK������h=ޘQP;�����7�Q<\�����K�U��7�>�2`SYe�,Y��|#��[v��V4qXOW����j���0�k�������Ґ�
ra��2����|L�0��|{���=*	~�r��v�$;y�|x7��KA�~9�W$�?"��?B��b>˿�����z���։�]�a�^�W��ž�Vgp��H_c��[A����?l�N��M"��d��ND:A�JS����z����"+F����hJ��{��+[��:HM�ĈS��p�C\*�r��,�ZԠF����cA�|y�Z�'�V~��&��l!PK�@���P33+R�Y#�8r�ӊQz��-]��� o��1��������Ld����^����,<�l mYv�-=ȥ��)~���Z����+$3485���x�Kk�_V���f��5O^J������A>����g`O�`��g�NT&�5�V���\�+&�z�#� �s�����١����w)�2�5Xi�����k=��O��?���AU�f���z��ޫ��L�N�'������b��]��q��ঃ[X���h�*��3-�f�QgE���|9�|��P[��R1í��v	(����Ȼ!U[�|HY�ô�dl#Ҙ�^��_��Io] ��t{�F��׎N,QG��d۬!9*fk�����n����1�ݦF{�;-��m�ւ ��M�"�(%�%-%�A�[n�L��-�w�%�5�L�dxr5+�˫��T�O�mQ�`�7�xb_�z���-�0��DL���Ъ�G��uE>$=����L��6��W�֌!J ��Q�ɥ�t/�Ù�t������Z6�)&Y+�E�z�.�l�&�qA����%�Д�# ^$�c@-��
�𵜗ZG�!YԴS_768��\,�.��u^@���Q����9������.w��&��։� K�)Se8O��[�`_Az�s�[5��y'�'s.�zSi_���S;>ǰ�>����^b��z#���፣�ה�V�" f�r��ڨ3 �|�9�5���ʫ�9�-�zqK|u7��'̤c��i���V�ϐ�����ü����n�P����<�-ߊA�,@�GX�BxQr�zg���vО�"�$�x�)��')�i��Og:����o��b����;�=��e����3�ɩ�.���gAd ��iJ�g�_��I\�d!�5`B�����}E"�#��
�K]v�(gc��u���@ډ]]�u�U^��}�u�b��/��f0b�ǣ�rA�Vn)nP3��eQL�G���?���ѧ}�G�9�r����	}��O�=V&��$�i�J�^r�Zφk�'�g��߫z��v_g�����${�b2p3Z���.��u��k��~Ӆ�OU2S����R��X��̵L�c�@}>5�6�����ģ�͚��e7?�
���\M�辰^��?��	�	6r��Z�RS�R��6��y�{�x6�E���*�8cYe9��%��8�U𤌥��x4s�+B)^�^2���,Vu���%����(-��BS�x*�Q��f,>H�&��<�����	N������(t&�iտ�O>�^1��M^N��WK��T+M��Q��~�:�#ِ��1,�³�J���Hy�Z�.��&�1���5��M]��h ������d�6LET,�Y���i�&DVr�}�K&�u�[�?��Y:���}��P�KR���D ��Et���)�5���k}�i�#(���Nt��-Gۡ�����f�D̍��Op�u�zL�"����p�&M�D�>��k|�/
��S�Π8�|�U�a�^|�Lj<1�Q����$�O]�	5Ѡ���[&,Q�1��jo^��`���|K�i&��z+��E�e$wa~���6-��!(j����vL��������*@� ����x�w]G.��G_���)L�(�.�P�U���D�����	K�%�x �m����ؚ�{���V�����dM�ʽ��d��o��v�R'���^+k�<搜������'S� %�V=g"�X����%{��2���Q0kK{5{��%R�Fc��oƦ�,ݬ������a��sUmU3�m��4^��x0��(���JQ
�3�-��B���Ѣ@'A��݉?ZKj��S8�$iu�
p�p�|	��R"��P�Ek(c(�)�������:�f�!�C��#85в����Zu�<2� &V� g���3@7F.JQ�*B�%�5e�+�~o{Y�_|�Z��[�,o���r�Ɯ�<�@�u.q�JotmT�_��$�Q�������&�p<�{�o�X�#������D�o ��,㳊o����Vʬ�Q(�(b���,�.�KIY���4<<�A�Xқg������d�M\ջ����<���=X��DY�����	�]���zO�}��N=�U��j����c�~�����e7�s��Z�ȼͥ����Se�p6q���\������*_o_x��wT�`7�0.�Mȃ"|�W��Y�#��/P�����y�Uỏ6\Rp�<�ro�Q*�,��5�%/���>2��>�EpPo�3����~*�1,���wK��b���S���=];��h^�<��]��������t�|�|�08q��hz/g����O�uV�aD�P����I�j$�������-#}#��8��q?<�l;]s�ynu����V�Y$�f��-N���Ꮔn���0��A�H�V�O��@�yw��:]*1����7��DP��
��6����<w�M���؅k�M������{��
�
3�7���i�D�ɫaYk#�Qq��R�ʨ���3�>}z}�ڎٓ¶y��(�|#>ĩ����S��6*-�D腖����M(��%�|���7g�=�Q�����Ǚ����>+�VVׁ���l>��}��ͅZ&頪-�,����V]e��pb'�M��͛g"�R�� ����.�lt~���Qw�2]��'��z��*�"��C{�:	����"(��bqح��������IY���g�Q���O��ɪn��>&��2"��	K�������n�,��4Y��drݶ�·i茊DW�ds��[ -�8VV˨�RK�w�!��S�M����m�2�v�nYbk��)�oD�����zm���z\���sp�F�~�)�Y�D���U�#O~��ȧ׮�3�N$�6;�2F횷�܌��ny����XQ���#V�84Y�S�Ǉ�Ĝ�S���m	�~�,,,._~��{��{>&.))��y26��=�Eb�e�����?�C�E1�#��ٳ>|�`E�+�����P�g�� `�����d��%���pFI��C���X�x�-mjjw�yP}�3���C+f�^w�V�c[c__�2������eͤ�}s2�p�ڪ41sfqޘk�ZL���]�u^�i�n�%��1��������q)��|�u��F��SB8���c5t�ʳ�%<2r������le�Ψ��jW�,'��Ix�Z�l�Mg��g?�y���ݩQ���u�a�%(�GF����G`R�E�};j����|��Y�!1�a�r��MF�Z�5I�� h0��Sl˞*f���������m�A�+e���T��n��t%��l.W���ׯŝ~��f:e�d���璤�����^���c-�:��|[�H����a9G�u]���t�
`&t(cU���`�H+^ ��@��l���n���nXu#�j�-�5MP��֫p�T�*���b��rCΌ[�d�ے&5-ms�Ϟ����X\6��Dk����˗mJ�&\�'\��~�|�&�+eV�,ɋ��:��g��|��g��k{Povk���}�2���.+�tٚ&�tQ��>r_5q!q}!�Q�A��ܳ�y8�9tu����i/짐�[��%��+�l�a(];-�J1�׺���D�h-w���ήO�����C<R68$d���z�y���/�̝��:��������x�l ����mjb�:;�o��ywo�`�a�ݛ2���⾻Nlw��:[0'bᑱp	�|\jj���F�Z�����#8�4GM��������28�35�(rx_�
g����bnS2��Q��/��U��%�<���Q�ZK�֘�8v�/�����w�|�k�~w�&"� �[�8���\� ��ML�_333wף�l����#��:Y���հ���Q����CE�.v5�!��9�'
***�ʞmb��Cf|��N+D�IXY�S9��O�KIn��]�8��Yr��k� U����i�F��wz��\�����O���@ږ8O�w_�>�B�F��VmlkS�;R���R�C>�\?��VY�s %�S�1�_�q��@:77gAh��@
�]G��t��F��FZ�����ugH���w��@*����ۇ}e�3Ma���fX�������6>t#���ٳZZZ�����"K5ٛ׮]�k_YYY&BQuSkVF3w�o��Gdđ��T^��- (P��AM��P9��/ ��ק	A(f�����%��-!��S�	y�*-�S"�,�<����,�W=%�M��s�����	2�G�i睕'��@�&K����&t	�38L��������Qw��Eo܀���/kW҃4��7��ث"l�*>�n҄!�� "������Mg[�ZJlM���^�O�M�ջ'��ӣx� �)���^;Q1�+W��ܦ�V� ���x���`���-�kf?�1��$Y�{lu��-�������a������kU��*|���:8zX��EZ-�)�\��+�l��Y(���3(Py�SU��~0���yVc`�D�w���#ώJ�=�k%�K�`�i�`��(�����ۛ�h2�r��O�������G���`:�I�b �WVVn�74�OAQ��Ύ�������[����.��ϟ_�����^&�(!�t �� 8�-YYN�w�-�t�47��������Z�q� �jj-��ROAw5v����YX\4��X��edd�.-�c!;00p���qe���S�'>Qc��#���@��/���X {M����B�]� O�W���Y'UŀПA�Xi���iC��߀t��G=V`�}�,�Y���|{��ļ�z�g����?{ju7H�3b!k}�O���;������׈*:�pv)��Z[	�߼k���%�̻x��sO�8���`j%�#yQ.l����	���ȸu�[������tmަ�����U����j�U)�|](2`�

�X�%���G�?8�4�B������S�P���zo��|xJ�%�` ��� �A�B__��wC�o�S���--��YBT�b<6%,@^)S�n����n���Pų�����h8���'����܄���A�ׯ_�����w������(d��z��>� �B��T�,����:Rb��Mry��e`��>	x��$���>�������\�ý�#̠���;-/���Z ��o@F@���ppqqi�W�[�ϧ:,#�3>>>.99BՏ�:�ֱ��2Vb�=q[Z��?H�*ɩ�$x����bC�f[>��������(�C8<$%2����g&t.,E������j�4_GOn�X���;c{>��9¡\�K�A�ҟ�i���X"��}D���� ӏRc:���M#����N�|�s,��1����ͻw��RRH=<`��c%q��o��
��f���e�{����l���%��}�!���|�;���pI���J�f��p�� �k A�y�N�������� �Y/��I �QGL��f3q�e�r
p�9k#�&`����k+�5�b��ٕ�m���c�^���m0ǇRR�6Rwy�&�t|u��ӏ+�>�3H��Sb�с�g��=j����������p�L��<4XB�oA���*��1��x�� P�[��,/_�\o�_��_o�1A��3b��̨ٔ��d�5�l��H>fO7@�ɩ��� k��f�.7\`�В�����1t��Q��5��Z��tݙ���¯_�.�4h���%$�x��1ϒ����ʲ�[���٨���߿C<��~F��m��rQev��R��I�Z�-~Q�2��X��ˀy>����o"�Tl?��^v��*��Z<�*"��kjz�v�IT�)(&����r's��z�.���B���K���%�c�z��.p�tJ��� t݀��Z>��h����'0���dN�kfh�Nn�m`����U�YYY�@���gL:�ip�+e�ˠ��x�����r�~`t9�����6�W��5�����,���*�x�.X�����]��sB��k)2��ǿ��eS���M+?��K�_�|���x�!��`�疻���\���Z>F�a>���:X�4t�IMy�ԋ!)��tu&��=.Z�MN�6�yƫ��g�	�	���Eؓvir�M�dC�ogK|j*���*-���=�N!S�q��_�}�be���k�J6��_|<�_�w}�n�˺o�ٵ��GEA���M�=���al�5�����1�~F��%�TRg���QN��F�3`j�IXJ��5�,��M)K�Vk��S���V�,�kų�B��]!�����\E��u-�����Vs�v���4�z�*�?L���T3:*�ZL���}������#��0h��Ѽ���u9]j0¡f|8B>�=>��llhʑ��R+H�^դ��n�*"�ɸ���m"���KCH�Z"tЈ鳆�!����R(��i#J�"*��z������)�Sn�?9 �Lz{=�4[��H�vx���t�;�/��4�^y�
v����ʢ�:�>$R�sI�����rE��ry|��kG��(�5Dv�VM'�<clЮ]�rk�U�J�W�)�����pҨ)���{��,��.�;,��hg0�Ց�Ю`0t�5���� �")�����%�dQx��)/Ϩaj��(0�@�a���hR7:	D�&f�R)#��<k��($�<� ����P��`='�����ރ����B���V?��P�.�Np�{^��K%�9ߢ�U���\��a:u@�v8�xP����1k_��-J���=C���t
����ѭ]����O��~������$��1��������
�Mo�����$N�V��Q�`���+��������.
.|��.m|m{t��d:_��}(�:+1��Bh��|@)�}��ϭj��+����G�8��F1� �$6�7�V|�~\�w�����;��l�'��+T�mOChMW�xe�}/�+$�+Xܒ���X���-����+�e���8!*5�s��OH�pA�O�צzoT���&WO��b��,M��^�YY�d^t��Mɖx1��s�-��R��O���%�|�z���?�Č�����x��N��Ô���k�
34��?u�cb���hG#ْw�J��q��l[YlE
@�_}��T��rjb��/��E�䊾��Jz��N�}N�u(M/7xo�%�D���Gkzy���Q����.��'�����O(���	<�I�_^�zYf0n��	^��a��5.�>�%G����u������{��/�+�%
=��tP#�ل�Q���FgZɀ�?i��)���p��1��_	�i���n�UOB��Gn3��"<��8{��?ޢ��0u܍+���&����:]7=ê�o��ײZ����'/i�*�&7�А|�ve��T��SR
1��f1�Y67X��� �gK�MbO J"N��Z��lFg��7�;̋��{��oZe�[��%�Z�W]w�ry-�E��Tt���|��g��(+%��mVF�r���V
`���F!���{��t���1�#f�:�}� �Mb��=	{�����ҏ�4�GZ(ٌ�c�]�S�v��a����2�o�Y0?j���[&3[(U?��ٝ��|֚��S,�Nވ*�)�w��k���ځ_��;�P��R�_�����ڥ��\=��۴�h���-��Y06����Jgx�eo���V��	>X=���1tЄ�ui��2H@h�O���{���\q����?~�osg��/?�MR"nm��#�wv��z��9>�Pb�ܻC�#���O�sl�V���;�N��=ZR��:��Б�5�5��%H#S���Y���ԈJ�*�[�5�S�;_<Y���Zz8c�Z�"d61:*�~H���.�����e���xD�2֌.p5L����0,Af��a��M����鉛�M��9'����t:T#�4�O�1�Τ��~Z*JE_�3�O��gK,3�E&Uw�!Mxf��<ig弝kd�pG<�o.�N/�f�rM�Yv�"���o�4�J�a҂b���Bin�_6���lNf��Y�@66�9[��}O�{��N�`�m��y��5x@�e�v�A���&c��b)OUq^v?9��^U�g�ev<z�)��Τl"���}����Q}g�c���<Kr���m�[R��_]�U6S|I��pI=�G+z�d���M���0���2��\���R#�~I�c��n�.���k��O��W
����l�	�x�H� [�|�d�-��G�)���|���XG�m�����`��xY-�ΩW>����|L��?ó��j��x��hwu�j��T|���k6�cwU����P������'$Z⋓D�GǸ�N=أ��w�]����/E��]�A�a,��b��Kzx�'n��I=A�K�����m���f*V��94��_Y�Yg� �	�0�5�}��x��٫T�ܹ_�ψ�s��#�:6�E8�ȡ.����uٔ��Qs%O�܉��Lj�un
���Ϛ�F�"���<k��#�$<�e�_�c;�Ϥ{S�]��B���*�G�7%�"�����
1Ѹh�74�����A�]�5�Fn����a���:W��ҭ���S`~�ǮX�Z��Q�:��?�X^L����츌T_�ܢk*�!
Uf�|1�c���K�2�ىy���gm��c�VO��AES�^tb���U��+zW�ve�r�FW��duOetL1�ǂR��	���q����P6g�oX䀱	�`�\�@�+s�Z|�l��Z��*_`	_���l*͎ S娺��v��L�e�'���27H񫜞�5�>m>t���8�bt�lAǁ��ӕGe��6�>�Td�U��v5�V&W���[��u���T�f�BS7�|�]����P!���i`+XzB���˭�˓d���*�6c����}]���?�[��,7�nN
X��o��j��hw��g�P�s���՚j~������iL��0�E��·�?Z�`��S�R����Y�G���yMg�w�v��v����QJ{��uﾛ3k�ڭ_m$|�E��f���>�K?>�ni�3���W#�ۏ���������#���Y9ϰ����)�������������mT%�ޤOm�Z��Ҧ�����1�$����e��������OD9�S������&a�5�|��~�+�16M+���4S��Q�Ta�P�Ż�5T�0Uf�"���Z�����^W\��&i���'���GHּ널ʁ��Zw������[u�߇���ۂ6m9�<|�5T��BaM�x��U����͝��LB��\��=�FN����	8�\�1v��)Oj���~&_�J/[ ���r.G�d�b�cb(��"�Z���ƗЊ�`�> ��{:�Q�: �p_޿����=�>�@�|n�A����_f����Q��7w�C]ڙ�{���l���I�=��>(ʪ���𲔿h�L2�tZ�/gޓH�M}�Srӿ�T|��{�,����SMށB�O#D
v���6��W�dal���}�-���.�27����������Z�S��!�|�,��u�5����lN��ᛶ���a�<7���<��s�f�h�8��P�9������IU�Ә�6YU�_����4Z��2Ѓ�!�t&��}�f��׼Hǽ��~��"�l�_c/�\w`���U���KA�ny�~W;�=�4b����{�A��mп�8'�Ge[�A�'����448p�9k����2i�%G��DV�ײJ@�Q$}�H��励�����U�Q7Ҕsy�Vp.���u�Q�ʫۧ����F�M\�7rО����Դk��>ω,�?��{&������<&��9:�l��P~z��z�#�V�'�E�}���O�v";h=7�r��҄��Vn����J훒��U^��w?�A	��	&1��o�v�	X.p�y�H"�����&�.��ɦ��}���˦~�TUF��g�U�i�-u ^�#o�N���\�V>
|��7s�bPσ�t|o�8�ԯ�&�ӷ�Q&mL����ԏJP�:�!�>�>��i���̋=�����2��k�l�I���	-O?�HX�����w���T^O1d�ר|������&h1��"��}����S
�=�?l�@�谵���d��Y�}va�����"�w�|�-�=x�gIY����/��N7���Z�xQ�v�?o���O��Ӹ�ygZr�̕Ũ�j��*�J��nX΍�nL��5��1O;�BH�A��{������xa��:e�92���ߐ�c�u�M��TA���4�/��^�S8.�4G���ӓ�7���;���~5Rd-!����݊�֭xjG&�W�'NB�(�"c�����k�6NX�c�F�[t�h1�{�oMT���(e��V�;�������*1u'���uȢ2�y�h��>�v�G�d����E��j��e�I"31=�b�f��;s&a�e!t���[Fnα_&G���8��"����K��v]��#U�Y�Nv@gqI����-��	׾$T(M��-�	&���G�rE�Kۚ�r �4�WD�|���]�,�ņ{�)�M�q�^6��G�w��E�6�(�C�'�\}������rIv��O�nXݯ�Y��\r�������}�*����&M��H3zŸ!�����y�);��v�3�.�"o,�K ���^;� ����� 7��Ss�
��#�L�n�X8i���&M��V �XV�+�$��=����r1b�ZNn�\���u=�X���z�����(r�;�[�>�ܗ'��̟�[o,�G�>���֑��mn��������+í?��<v�ny���g����ӡT���O��sk�ϛ.4����vN-PK��d�d�|l��Ԝ$4.�P�3�1!�^�s�U�����`����l8�h;uPD	�w��.Pz3���}r���Tu�͝l�mEUZ?�6��Z'�|ʛ�x<��g��T�����g/�e��RH��(vt�a����*�(�:�����J�Y��[��v��6'"u���a���?��Bqm0E��,i��v~DnA�
��
@�=��ޚp�H�S�0�(�����t	��t6(�4�~la��V���h�mﺶ��+���l �gk�jX�*Bu-\2�k�k�_(��T��{��T��\���ȣ��9���e	����ҹɃ6�L޷t<�%�^e�z���H���ll���@J��8�v~?{�H�p���~i�E�l\_϶lVfv����|�&�S$�����K��P�wq�X�O��@�<���D���	��񕵇�O�3��}��r��)��i�t��L��7m�g��#Ο^~��v��.y�3��	�k�W�jj�?����#�����P��O뮥���1*{�.y�#��C�Y���j����LU,�1(��o�$��-*fiX*�����R��Ь��IN6������Ѕ~az���o�<�̞7l�2�[�qg�H��N��X%"��~��-N2q�&��{��!Di���C݃>ц��~�w�V�%��?q�i��2č$_�Z� @
cl�M�O����-hN��|M� �f�\
[����T���H��n]<OFV��k:&dQ7�����d4�lyr�� gBrb[t!VV<�n��LU-�� F39��C��nG� *����;�{��Bʠ+�xk9H�pڨ&|�K�Â����0k�&-��K
>�Y=����#1Ix�$�/����W~J�T���?��#&
7%����guЉ��~�����;�-c�.m�W�W:,�S�"�O��heY�}��ѝ�{|Ӣ�~ �o׷6X����{
�#�CZܖ��QM��%Gf��~<�X�\}M�O�]HM�Hp��m'�1m�/Yj��%?�6���][/ �?֊Z�=��2us��ʹ���̽r>�»N�7�D�u-���\��a���i;�p%�d�������5�W���u���uU�i�7U���t㳉��L}\���;��D��ҧ
�Dw���`�=	y��%Uٌ��c��\:h�ˇ,w��]�K)��-�]7����J����������>!K3;��Hu���v�1ǊyF��#����۞��o�IF&&I��͉���`�}�R�[n�-��%��;4y����l���"�*�傶�i؈���ƝIuz�����?�V%�.Q!���	0��ǨtͰ��=�0��@�k]���X�շ�E��ynR�w=f%�U�H��OkY�WcePZ�]�WtKed�׾�U�ǽ���)Z�#�-�H#ˮ�w��^x�߽s�����h�_��m�I����jD�����=C��}0��͕�/�1uX/n�$���⌥0yӆ�{�f"%�[[�+wZ@en��L�m�­m��T�	~�K�ܢU�z�G��N{z�kA��J���ػ5:o#����|�y�6��K�EW %�BqǇ��{H�Ȃ�>;����ҕ�2W	f�/J�p7ܤ?4G��c�4�Fݠ~���$��!N��舘�6:;�3#��(x]�7.�՘W�5+d�����n�s�L�}�♽��}�n+L��q���OPG� Ǿ�U�N�Eźt�E��I�΁�*:sx)#q�$V�8�Ö�?����T�F2iA��]�aXҳ���O����#�'A�a9���1h:�$�L5�M����W��=�uY��$Ұe����Gb7Adp��C"#�ʤ�Qӯ��r��ߩ����}==o=�S���*����5�~�kJ��	2�j�N��^F����x���%*��ˁ�ѰN��n���"�b��@�������
���p����ܸļJ��q쀠�\�p&$pڌf�7�_)p���t?���]��xb���b�����X�>W=�ѭ��6���쵍²hs��>W�o�ԥgs-c+�������c\��\S�V/��q�/^�|5�"�7���~>ʦ�F���"n��l�I���C�e<��j\�݋ikk4tt�^^���4?�?6�ε~`aeͭ*X=׃��̽�������AI{���^�����E�2���%�t������o�9G*��g�bX���C��[۽�E����o<�X�~������ 7U�A���d)̕��Ъ�f�[iBMPSc }�x�?��wN�l��K�N�Ol��t�UN������Y������	Գ]��9�/�췔AA3�M�&I=6��\�����*-�><r�X��E�����.UwOϲg_�N�k^~�~����o)~��O�	�ݝ]41��
����Z=�SYV���2j����D�ԓ���,_L�Dq�s���kF;&ƹ���׳����Bq�?���l�K�&��LϞ,���zg��=G��������C�I��C4@~yF��Ӎ1p���ZCo3���I��.�1o���7�7�+w�Ztn$Q�ˍyo�mPI��?:��tE;�
eMz?Qџak�\�C�)*���kY+��:��©�/��؞��()���l�ڢ��3�nL>��vU�-�ݫ��
�c��������\��?Ѷ��#��Q�/�ǣ����3�3��Fgm���گ� z���������W�;�SV۱�/IA�K��"�>�*���f�n��ճ�V��/����SC �Ѷ�r��.�Zq������Է�Q"�c�o��l�ݯ#�Z��we��4�����M�~�~O��JJ�#~��=�Qj��層7?2�u�x�����h�s�72��\[  �ہ ���@���
����:-���Ǿ���1t����M"�L�_����ݷ�<H���������gB����[��ѩ���ݯI�U���L2����4l�A{u��f(Ĝ��0y������H�lU�0�k羜��������G8s���/�%��?=���( �DII9V�ZYY9GK�:��Y^�3-ˍe/N���w6��Rgpq"����Rf+d����͎���q�Iu[��h���1A6�U�w��t�m�mI_�K�V���܇�KSt���Y��y���mɑ���6�8�F!vj�;���&Y����^�9�~�ǖ[ò�ي��,w6�b��v��\/���!�nPQ�&rQ(KC��R"��K�IF��q���y.��b>`����i
�D<C��Qgi�v�\��̊���)�)����ƫY�&(߽�>!���UI�d?l��/��F��*!�
�[�yz��G
.��"��޻��K�8z
�t۫�2~d�;#���W��_*��i��x^.)�{Ol���k��j�����f���aEqG9�燍��bl�vm���5�����|�ut�P]�/H��#Qʪ{��;��}r��F�V��
ldc��?��:V���ԮY����ٗ�6�3��L���dq�Sc1Rl��\���.֬��г��9�1w�RѬh�zA�����f,��N,M|��Vr�~����[=����织�6C*E��(T��W���~���Y��n���p���ۦ4`��0���;6Ϩ������,��z*�9H2�9������#�������x-�s���G2?�FY%{�����z��rF&&aQ�ku��${��w�����R>|���ÿ��Y����`?��.�	M�6&b�&�$��m�g��a����餽�Ż�����w�?�fx�9xh�VT���w%����!��[9>ݞ�g��=֞Hx�.�5M|S$ϰ����\�����b|����{({8/m���ݕr�m���@*쬀!�Q��� 7>�9������OC�6o�K*:�%oɘ䀵@&}�5m��I�O���0i4]��be��GQ��b�Z��9������@q�.�0	UN����t9�-���ChJD��9�;��������G`�U�ׯcުuO;,<��w������1`�Z(r,[����0���L���T�h���|�����fǅ�Մ�����=����,�t��>�e���C8'{_���/~�&���V����X L�'�Ĝ���2Qn�9[�~k�$⾇|d0�_h�-�S��uq� (mc�a�_:4���ӡ,Zbw��q����|;�\�gE�	��W�刲5�Z)������w%*܌'D�uVi���l70лg�+~���D��U*�k�s#�D�m5n8��t����b����b*�DZZ�[�0k�' �4���V7Y6�����թ��|"
�{ɩJi���Q���ꫣ�j��		I���.i����;.�! �� �������ݼ}�k�뷖�׽��ٳ�'f�:h���gA
!�`���`��ŮRϋ�B���?g^��:}Lv
����?׌�3�ٙ���ֱџт�jڸ�����x_6�	]���V}]A���Uq�S����s]�P���K�2�BK��*_����2�oi��2�g?��$r����&gf>��|�0_i�!*��0Ǯ>��ֽ}�@���=�o�^1�f�w9�˄��O�fۋ�4[E��	ʹ�#�J@�0>��]�t���x��:VHφeO�7=q-q�'n$uArGՠ�;�7��~gM�e\����&��A�l��*�[j�q7�[�7������@������> �&&&?���\\8m���aS��Oh*���-�;�}���ګLW�2���P&�>�MW�h��:����QHJJ�o����E��������`�T����pu�rf�Vw�%��cν�z�-n5Լ�>RqݗwDkU+��Α�m�
���+zp����E���-W�v�`���6NW�;)�;�6����o��i�z;���2��~"Q��_�	f8����Fs⨕���%r Q�jJe�%��+\���,��)�ٸ\Xn��Q�s�8u���P��/Fk$D��4�9~Q�f�Ka}�5��՛��L��S,X:c��u�~x-��fC�p�ч]VЩ�W��C�3@J���-#���/$�wv��&��<��)���'����Y�>��:-݅�ϝ�hr\�O��kʘ]$���]����`�[�-�,]�׷(� :������Nr=
�Vf����Z��Wu��8�#�H�(N���@�n�b��t��{f����'}7h 6.�~~(�v�H����B\wcy�ߺ�z����w�[��X���+Ot�K�m� ,֡�sY}�ZY`P���9��ZT?-��Dn��A��/�{Nl��E�=Ꝗ/���D���ޯH �qd��-1a}9��, e��.[�Z4��\Bȭm�"Y,[��8p�̫M8��k��x~�ҥ����t7U?Rk�,�NS���("*��0����f4���M�j��;_�V�blVR��J3c�l^���r�Q6��'�+hʘ���:��~Tu((���kso��{S�;G���c���<�Y���o�?-U�%\���&bшy��`p�
|)����\6��	�]��=���U�>�6ŵ͗N�+�u�	�x.MS�j�Qw^&�������#�	�C�$#q;?��IT�]׆- �����_to�6��|ut1��@ ��S8�b}�t�����	�UZ��s���l�~`#�q�v�iT8��v�J]�/��w�S]�s���ZE��/�A-���[��Z]�?[��n'�J1�[��$�U{�u�t��<l>�r����)N�E�1�-�"��j�����8${��k�w�c��~@�û�����f
������0266\�
}��F��F
��z�\r�;�_6����%{"Hf*G�����B�P:嬭KÉy����\�W\���x:�����.5��l+�KsѨ����8���9�'�rYF�)�qH�G�bG�Ƀ��N�s ��8�\�q\Z��,*�H�y��}�38[4�ߖ0g�	��ꪰ�Q��Y#55�)�L߳U[4�xj,[4N&����<w>�	Vl���¤�Xͷ�a���>B�r��ې�{<ջ�
`��-E��j2�ѱ��V��Y�6�,�Ie����h+���N��4o�\��(��4]{0�*M#~�Ҫ�g0>Ѣk���I#y�����I�E-Å�|����5��&\�u|
^����Z���4)���)7dI:B��@nב��x�����v5�ԫ�w2YB�~k��'z`GB@'&O���dZ�l���A],б����=��m]�@�f3+�f(!�a��){oϔs���
jA�%零6Ie���4oqNAm?욖#Z����@=s󺍈r����2��8<���ƌ�PKg��3Q=�s�da�.Oч��G���-؋�˙���vb`��6nX3d�E��M�pB�/��{��v�_����Z�$:���z
�c�k���Fprig�,o�'F�y(�y���O��¿�99�l-��>����Ikk�{��� [��ʲ��De&��u����r�e� ��ן�^vHrK���b���6]���2�+��~�I伤��|�bra�Ȁ��aX���1�Ԙ_M�
7���+�6�1\l����E��˓�P����&N��eDs�[�}BW!�z�a����[�y#�ks�|Ec��Ы�~(�j5��3�{�χ�gwx82M��/�@����<`
ŝp];-�<-�dQ���7��5�������ܶЯ���Fa��_ �oG�U�m�!Ł��:'���M�~���f(��2!ޱ����q����b��tQ�^F���+��U1j'J���:���q)(��;�� u傄ל���q��~���Ј�S�9'�iOV:i���p�}�>̌�:Z���h8n`,M���j���/v{ЛP8�͎�woT��1�o�("�#�6�t��Sj����x�� Iu��R!kwö�T�eU�.ai�g�r*�sr{��">W���j-?�睔E��������qnG�fwe�D��c�'���쏐+$�jP'��}k5U'M��9���f^���S� qS��	3����;�j����+P:�D�^N�3:O3 �ٷ�zi�����3�˴�p����#���&�γ�-P��xwO�UY���Ee/�)H��������j����~YdR�@�@����,"�C�+\6õ@
�ǉ��iz�:������?�ޔ^�}������y����o�w�!g�;�J�p����
�=���r�5��0�ζ,n����^��v���x��J��=��ы!g���@��c�Ȳ*].�CG�`XcLn�@ɸw��]V�T�i��zV�/1�='1��������/�	=�Hjh���|�7��`�s�ɂ�����N[cd�nksŨ#������[��A]W`c{�b6���QLA�Κ�W ��Ư!����\_��~�Wr6�X4o�������V�^*��s1�k]������]�` �b���U�b\�R�lU!]r^#������ےOn��7�^G��)wN�.�-:��"�*n=���Ϊ�}�ҹ�Ds�����e��y��z��5��'PP:a/Ԝ�RDu�[?W�Ν�v[b^�ѥ'�C�w�ާYo��Ov�*���>.�J�M�.i;|��賁�)����i��D��b9.5�����AY���
��a|	rX�&���`�rd
�NY��aW��x&v��e�����ӯk����t����f����H�y<���N~(����J7«���V}�l(j��@`���j����]o�R��h���d�6��ڪ��\G�� (ZaEQ���>[�V*��1!_��1Q,��Ղ���4�!s��,�D���X�QQ�c�Ub�a���~��,י���\�9,8��n�/�mfnIƠ������7?�[έ�o�nl��B�R�@��v	=K�7��2�L6#X��t����]�sX/[�_�::k��\�L��gc�P:�X����qy{��"DǺ^���Si�yH�!��r~�PN�GyX�?Ʀy>������zq~���sm!�o"Sn�;Ѽ9��N?�T�Y�ug��^M?�u�I�C�?��Ȓ_�@S`���G��>� �j��x%'��L۟b's�S��񊭙7��ːg�B��h�@��[�Y�]�,�Ѻwwq�i��b�$R}/�f)��H���)&�4O��i�Q��z�`͟��!�O�2���g@9�nFS�E����r%M����rK�qz�Z�T�f�µ�Wi �8��U ���E*Y*I���gG�!g
��`�+ege�rZ�l+�����Ub,�HT�����-������}9r��1G�L��qE�G_�N�6Z���;+{���Ji}=���?Ϥ�%���o�b�B���T�#��#-�E�v��uu�u��spqH�	$��]��M�����q̦g��΂~]9�BH3`����Ux�%�5c�G�w:��=^Y5[���Z[���e��jrj*���e��yn�T<��x���P���R���˕�����kI_��:��&:�[]	j~!k����yk��4 H)qpW!wkyj����-��-�����&NO$����"@������){1M�,���R̘>���q�`�I`��:��.�Wx��c�q#�;�����{��LvS�Ԋ;'[�͢*��X5�[���3����tb4�h9�ˌ�`X���;w��$��"0��UU�2�ܸ**�1,\��dW��<������sj2�gLlx u^����՞�c5���<.��[h[q�4�ܻ ���	�²���Z�f7WS��-v'q�"���sX�|}�@�>�dn.��jO�t����?L�DmE��>$c[b��@u	����5�����	&�38X��)�� �|ӹ��>wZ3T���O�*,I��jߵ���U?�~?���6ku^��6���w\��6�#K���O��v�p5h~�!�]�>��-�P��*N\�����xa`IjC���{qq��!߿$)��=�p6ǜ�����4;[�/]y���-Nˡ�@����<5���I�>�wW���ę�]�
k����������؃�b�G������4�a�έ��᠛`�.+{�c��ȝ�Ool�Y�M"�#�9s�e~
��m��T'�Ѐ�j�WT��.��)+G�����_a��OMMuU���k��Z��~j.�#���ƌ|=����J.��pX1~7��n�Ѝ;���#u򐕓
{\f�F {#D��U���hH�a�*�./��c�+�@�W���G`sZ|������ܺZR@@���{��îu�-|�P����h&X!�z�-�p�������-�pj�uۙ���D��C�z5�&dt��o��� ���,b�nF�љ-="8�D;���5��l��K���Г�]�0>{lI]�����'�i)s��/Јgl��}Ϡ��!�U��V���~i�p����q</���F���+^Qk���!m�+׏��2�;�t�� �ۊh>���i)�u�2rǻ,�/�2��b�m��5��m����e0܌������*��}��W�"�3��%`H��T��Ԍc��*�H�d�=7@4&f�4ܵ�;?�2X�^�P�1$TҒ�l��8) ��*U���\Ξz+���7�(f���JCe�4�&1.n��><.WmM��[��C�P���R7�(#�.�<�H�jW�I���r����M�B;[ۭl�RO��_�����s�w�	��Otn e�'N�w2&�����b�5��t\�������k���&g�1Kn��n"߭�& ��+��	���鍄����8�O��8��*��Z9М3��C�j����D3sM�������;����r��4]�l�����V�:2�����CrO5����Ԗ�%'ۏ�Ѻb`�]+,��OR����p\�2a��p�gXgpѴ$�7�2q@>�M���q�)~ugu+��d��=�K<V���[�쌅�9L!�)o����ɗ6��0�6�B���B��U�O%	Je���i.ogq}K<��@4d��vJd�o����K�������lD9����t���fb�B�S�8��oS�90X.�;�n�%�҆�7�o~!���h��o�\�-��Dٟ���ɜ�� ����:|�-g�k(���V�,.YȖ'�-��E���mY'mE�N��`�����z;���Fd����O�Q�vtg��7��ٿ7&*��*�r+-~���-��E� ۜ{�4�K�MD��W�r���_���x��$������N艣�B	$vk6��Vv,���1��j����FQ�vśۜV��&�����}�J?B�����dI!a���+�x���Bf�p���;���o��ߏ��&�m��'�a--�BAw8�[��D�A��:7e�u���'=t���a��Y')0л����� rͧ�;W�q��L��٠���5�2���­�ŪϨwI���6��>Ұ
U�z�+�v������#8n�o�۹�&π���D��� �N��q荩�6�71H_�����u��Y�_(C(�����/��̠���ߵ��{ ^`�\OZș�|���*�{\�.��ذ�J���x�s��ې39�Z KS�8�q��el�l;"���_��؆��>�:�0�Q���w'�C�;*�r0��_cF��Ӷ��H�ݟ4��+þ��`�ۭи����3R��e���}60%�2=��-�U@��Bhf��RvXeN��[�h� S���?��������60��&�ч���(��4�M�A:r�ŷa��9
���������,(���c���3�����3�|�,��чno��ԣ"\�{��d�+�/C�������l����������RX�n<�a�&�����Wqw�d��]�RrHv7`0���ZV���MUT�E��� ������t]2�0|EY�[�r�@?�4�]���*��(,�')��h����ۣ����f?Q��[��E%N��W��K��^��fF 'c����%����z�c�ß�׼;�h�����*���r�.�Z�1B�֫�&�ޮ|7�E�!
�A��AE,�?��n�B��P����V�q8z1"�~��冶�.ɥ�_W"9�#C�Jo�[өܘy�,LF�jucs��K*��lp�u�d�6�n�t3��6��|�wc��$���Q�5T�4s��7@#��P̸�hr޹m�����$y�4$�r'���*;bVnT�#6�|�7Zx��l��\A3�/�灊7Hf|��������U�8o�����Op�,9.H��n).��{3f�ƫ:h�PV�M����q\��b�U�p�/�lo��P��8	+�^-WߣL�~��t�!z)&�^N��˭wԾ�[�)���X#��_�B�m�:�&X�o�r�I=��}2ǧމ��lor�����NB�s�{#݇u+��E��������;	�
�U�����2�dFVݸ�R<�x��=M��m�1�)�{ʏ
t�㆔��h8��D�NJ���1V�(�߹�����>;�����h_T9{L]��"���BR�����3�vBNQ����q��h0����d�\��W����G�I�� '�b�9q�yk��5�_��|��~�T]�~�x�Ҁ�gb�l=�k_���-@����"VX�3���z�����D�#&���h�jY*B�Ġ%�	?�E��j@O�h?ǚ��8���m�`6�l`@�͡B�+�}�����<���f�Ƿ�t��kv4��A�h�H�������v�?
���6i.��Z(�K��.^P�B�������qC����=p$��|*���6/��y^Dx�ݍ��/���<� �t�߻7�Tk~�l���F�b�����#:ZE�x\Z��<	!���p0Cᮉ?xG��&.�[k����#y�g��?�hv��.bt&��S��̱@ƣ��ׂ�,R�S\�|X�7��W�G8?�P��e�:�����ƹ�̪Q��2��O̻&����q�(�gR�x�~�O�A&/�#�����s�-?s�p�F`䒘�p������:��=�?�Bvw=q�[ȗ&8�LY��y��f������Og=5�U�6Uv�h��6�7>��*�
��
F�����I��v'�i��twxB�v�V,�+�7&K���t�*P�NQ���k �W�u�DW���C63�EVȄ.W|���DX���_��h��H�x�f@#o�|Z]=�u6��A��H�?��|������89�Y+X�B�X~���0��V+���ri �rI�3�Rc�u����������$��Ƽ�Ƶ�$�v	C-r�+~3!���@[.�.��a�%��4��/p��;T%�::��fO�	�\x^�� >�ccF����@D���s��d�,����d�V��$�(#vu}i�)�E)��}�*PdL��~*����{-���Ћ��s������������a7����,gT@���<a��i�R_�l���R{s��#sM���t�8\0���0��1n;s𘯂W�d~�Y*_y^�
�6�YB��vnk�R/2��"d�P��7��ė�Y�S!�b���M��=P��|[}t&`��L*�ꚭ���	q(&Q�����d��]{�PB�U7�*��,��0O�{%s6�c�$	)K����B��RfGĂ�>�JG)^�b�������g�V�w��yA�_��(�=���\�t��Yz ��g�	������t����������N�/jZ �	끏!�X`��e{&���v<J�"Ll'�R�����>����X�G^�}����/L�`��xV��D��}�iWہ����5�E�GJ.$����zݔipܥ���h5��D�ap[\c9M���ao;�X��8�f���M��O �f�=U�U޽~Vʑ�cO�</2���)��_�h�uH�8*�	�R����/ރnd�*+�O�-��uoe�{� D���(��f��E���q�;r�uFJnL1A��-\0K^Z����\�����ܲ]�fނ��6����/u��D�uʦ��&]�ı�W��1i|���2�e���!Ce�a<��r:����ѝW~�ں���b��.��3dk7�6Ey��p2��=��I*�p/ ���A�k��v����??�ϴ����;�F8R�2�hh�e�>��6�����GbCfG.�B��Q��d67�	˃�Q!)�,�
N�EV�������UxRDS/���x9I;~������-Lp��4x^b���ʾ� Z(4(���Q��!�d�Ӑ�č���gꃖ���/��9M�޳���uq@��G̉ c"���/R_�X� �q��B.�_�-��^�.��v�1��:�˃�T]X�qd��Z�z�����,�~�adpz��\6��Z��t?[�k���t�y�c7�Y[��)�}�1��w�;��7DKA݆�,f�Կ{"��p��:I����U�2��s0"�Ieg���7�#[���e��'��9-՛�ff;����Ž��D�����@HÚ�,��\�������MB��%�$��y��jah�� M�*�]�g#F��n��ם�RSfr!��x\�R�ֶS9���6J@�x�^�^=s��_Px���l���8�7X#����~m�E���}�cM���������]W���k��Qw�5">I�d����VQ���t2y�U����8foC��s��XV���%����	��a4-?0������a���R�F�֍���ϊ�O>,:.�Z7c�\%��oA�<\X	��Ko��F����9B�/�!���`�x놾|�R�/S(D5����m]�&辮3l��Ê,"A�pT��zOoqTs���� v�#�(�i\� ��q@=8
��+S��K{x����g��1�����ѫhN�2�$
��ݝF���D@�m+8���nZ��R�4��-����w��Z�ۯ�g`�y�:Js/w��rdlUW���L�C�t���z�=�w� �"�z@� C'��r��&"�'wd9�H�t���V��%�bK��D�d�$���%d�̄LqNE�����(�����8��l�Ƌ������;���n}��[Ԏ\�֟A�YϬ�>�#&v�:�K-�T7��5�#�<�7�Y������-Da>����xW�j����ռ54��3'~�3��nf�
���M�����?|��r5P���;Mس��k��ȿ����HD�?y��?����v���J�� �
F;�0�������=�u��k,6�^�c��" 
o�L�=~$�5��Cp�g�-0��M�ScW"<?�ǧl8�r��G��Jm䏵_ܶ�l�v<O�$��s�(�_Ĵ6��&�@Q"xB灈Q�^&Ic{"ފ쩻>�1[�c����]�x����y�x��앐�����'l�~��6 ���R���\wT,�>s��h�w��&������$�tG��� ��1g�]�����6�����t��� ?�ґZ�4�W��_�b��L�7x.�O��H� B\�AO�k'��e ��� ���h{��6�<��L�F��2�oA�l�/O����64��&,<;���<a���!IW��Jҧ)^��h���5~��{��4p`���VgV=�����N�dc�K�#huP֬�f�3v7�C�Ж�>�6�;�ZE���q��\��v����
�ۮ՜��[}��?�\� ����,_���٬'����O�5��ϭpd=Gu�t."ʌ�+i�|�o����g�`�O����%f�W���She9"�yn�����t������5|�M�����B4xY��)L�ؕ��ytA��������0��`��\��r@�Yq�Q��0�lg<�Wp?��Γ��pj2�E���G�x��'�܂��<�t�ur�=��i�Q!fd��xiF�/P��K<xV[��:<�j����Y�qס�r�D|�u�򌘝�g�
(-��w���#����[	���S�V�����|z(��~����O8��Ĝ�[��@���&��eґ���*��s�F^+�Ӆ���9,��� ��������v%��ddlŠ�V|�K��8���4�.�Y��&�E3켻�`��La�9pDtj*f��@����]��0i~�T�L��ޢ=Q����C����tq�誵�u��Ċf|���͊���&A��|b�哺�t��v�����MM��V�ha`!kղ���t��}~se|�o��>A�/���Ć�e^xX9���3Zi�z.�Bw��_W"���;f��3�w��s��'��~Y���j�ʎ�yw<�	{}0R0�Z���҄=����'f�����M��9�װ u�;�������?�5<�*���	�4�!�d��{�}j=�daQ�ڢ;�k�7��M�.]1�-O����?�H�@�����y�${�Ǭ�0q�4Yq/�6�,o�>!hE�Y7?MCt�h&'������hD��1_r���T���L�y@delI��*�9 �4�v�3��LU�@D�d��9T��p�/S�H��fn�.·\�M:�M�/�g����É�pY�]���S�s�l{�㢥��e3㇔�#q�[E�ޢ2w��U�	�c�x8R��X�6�~`Ϯ;F��������B��	�g~�)|�q����B�)<!G�zO�L&A5ے+E����@�9�	?��j|cr]'p�e���^�6����?�Q0��+4��-h%�O\�sn����0�=���	!b�"
|�$�'�noMD\�0��ZJ�mUW��Y��)N�a( �7��_�!o�]���N�>��J�����򜌂���W�d��$��d���Ό����P̘�AQܸSV?߿@-(��_"��=�yP�Ϊ�~�?�/[�H �Ԟ��~�E�'2��l���}[�[^p��`�q�w�ϕT�6�WG��ס�
�{���0Gx�]���s����n�5�X`xl�>T� W�S����7pl�!j�.�þ<,�7�G~������i���s���P��Z
��7hF�Q�ǝ����*f#݃��m�#5�k^��2��qӟ��7g��R�K��ϳ]�ݖ���ի���oF��:9h��v�~~��OZ8<�U��LJ�*A+&v�����Z5���?�yt�&	9H�[?[sX/�M�\�D�e����+�}��#�ε�v�a�w�"��%���$Wݮ>�������k�{�����+�P�ho��`1��s�Ցl�}E�?��X��5�i�Jn��;|`]����ޝ��Q����L�4[]}=���.G���aݭU���oI�I�N����{[�el����E=�MX��O���8���j?�[�乏`/�����X~��������^O�^�]w��s�?����ZY�e��>5
ɣ�r�$T@2&Kk)�����N\�O�a������pM�0�~%A��v��9VA�Ŧ�!�S�Uޏ#��O�0B�J�PPB�_T���"��I�����<��y$�oXʟ�<��  L���6N0���w�֟����Y�o�l���G����V���«��v`�Lxg�Z�&��`B
�-�nI�F����**6��g�VH:l���Hx�a&�E�|�nC'}&̼�|�&�וt@��7���"�"�)��#�y����Ñ;I`�4g����=�$�*�&�MP"����a�zř�h��}/�o�Z�H�̓���[m~�y:0�j�L^�>�˅�."s����+��������;��nA�`�|��c�]=���O�ozY�:w��It�R�ñF���eK�!i�*�4i5.�26y=�uJo���-Ԍ��΂���h�&g�`��	u���?��g��ld�,^_�zrOk����j�*&���
i���1\�mE����nd�*�;�:�d���-�$�a�.['ܲ��Qj�cX4�C�~3&���?�аdx�J<a�Z_�?����O�HCi�^~<��~~=�]*����?�Vҫxf ʑ�,�)�R��	$�b<:��:$��Q��ep"h�s��
��bo���ǛJN5]��{co�^�р��;!]:IO�ig�`d
`�#'R�/7&[@��#�N�J~�t���&�u@=}YV�#��0��s`Bu�?8(��ƅ�A5Q���q�|��C��|u T�kDx�٦��a+d�;7���H��fBxT�=�)c;�׺��'����S�>B��Tc��������+b{6�*|���:���")R���5�o�*ctӡ�����,X�WgXBVb=�5WX���j���#ï�rv���B�@���IW�w�9R��&%g�,3�K�Z�QL�=�>��Aw粚��Hi�\�����[�����7��q��)������Oo~=���m�hF��>�� ���;�p��0�$�a�K�?Ӈ�.��n��ot��_N���x||��	9�L��eU��;	�ۀo4a-oGAh�pĵ��_�	�}���zLYPPho��^c��"�NIP���1Q�y�t����F�n>~�V�^��4#���B���r����?AeWg^��[9�Ђ4?�'#p�zDx�D�9� �I���{Rl��dw��Ikn}JA�kRfܡ���#5�I�v�?z�z̫�x�;�?�%��*	D�]�^���� U2��RX{S;�m����G�gS㊄�����}������@:�nn@斫�c�/b�c�����t9�ޣ���>�I��f�6������21����'����L�Q,T��{�p��4�n�/�QWX_�ݱ;�
:�_�'B6��u��)Ph(:H��~᝽(�(�,z[���˲?���dt|P����й�0?��A!�HŖjHI��d��E������m�cl?]X<R�':�:A���1�f6Z[���29�|�*������P��ܩ>���#
�y��KŨ\�["��_�w����� i�fU����M���vj��$��^xԪ�obc��A("��$����E[)�9�4<cX�gs���C��!���_��	�����0vA�4����br����V��V6 B`�Lǁ���'�,�7f�4��S��x"D��"�W��m���Iʾ��]�u��#�![�_�~��gY�$���Xyǃ�YpP��������E"���6S�M����e�#��=���W�[J(�Sd�9��L��`L��<;��ʡm�\��`3�s�
�}q�*:�@YnU����QTY҂�Lγ�{܀ʅ�a���?�)߮x.݇н�K�N>	� �����T5y�O���ݛ�#���&_��*Ţ��4�ն�3;|���#�A���w�WQ�g��X�A2�����;�}�[�����ăV���7�܍t*�����6��+-��N(�=�)9
=Zcc%e^s�x��]� ��6��6>g�����f���4A�9&�b���K��L2��H0+Zª�,,�f��;�^�k��*oM����p��T�9&|;z��2�Y�Z�H��z�ƞ��A|��s�&+Wh]Gk�Ll'E.5��]�-��yYn���30FV�̶�
2���C�F�]"zk����<������s����غu����~It�C�'@2AMU>xO��1_|�:-P�i�f����mp�1�ɂ$zr/���P��C
�jK�s�lvOk��y+�ۛÅ��ov�RROo�O?��p?.�֯����]��ȯ\����'��5y���G���Yuyͮ�.?U+~8�&��+��1�V�>�㜟j%�d�I�G�Ǽ��c��Z�rXN���R�K�aN���5⿫20Q���*��P �	��|�ł��������R�ό���W����|j2<�I� !-�f�ܧ��B�g5��^guz U�N3ڈ�	�f@�U�@pz��<w%������~p�@4�(�GW9���8G6�_�A�p!�w�)Oi.���u����������jn*�(��= ��n�٪��N��f�Ґ�Zq&'�����!�vez�4��|�}��"�شݱa�R�I�����t�d����a�ΣR�Ƥ�����-G�������m�^|�C�i�G蓲���o'U0�y�>��}}����.~ُ`�8� %<ᝃ���ҏ���HR<.�/v�G{t��h#�b5P
Q��2�"�7_�! !�IG�
���+�w�<�V������}P��yr;r��3^o���Y
ْ4�Jj�x�t�i��؍���e7��X��?o���F�Oc,�v�I^qG1QY���f�m����V
�x�:X����5y�_��P>5^<��7u�|�4�CK�ɍ�}�Ȝ踉�<P)>�̘i�Sã���y��o��.���S��e��<֍�j�խ�-�eQUb�p=��&MҔ�^��⥽r��m�
:P!Z��8Q��>j���I9dX$��HY�A戕(>��_D��sAt5:bۆZ=)�1$���
T0Z����l��>?�I17�itE� ���sE�RZ.G�Vy�j<��`c6���f���XX��֫��4���e����ӵ����\�U\����[���1�����n����n�X���G6�l��]2o?�d)�doUǔ_ ���Jc���.��I+HLG'���:Pά;с�)OVGwm�!�۝�N���!�v��d�	}�Ӽ���+�)���`�<Rn�h��}�Z��{��0�/k�b���2�\��5�xk�.�ϵ�B�c�U'��tyaά������g�@���z��C��5�ڱ��16��C�2�G@����ߙ�E?0��������$�U
����I�fR�����<;)x�iEV�@Z��kZ��@=M;�Bw(�A!Q�AQp�N�sz2ɇۉ�'���|����nB�[�Ah�#J��L�����
�7R	����L�ȅ�D��ޛ^s&�5���J������`�M�������M��i�g�x�=��<�ț��t�|uW/��w�K4D�F�D�־���̐�W_��;��M���s���-�!�F�[?#��]���9���g�d���ȿr��m{i�Y.��T�����|�Z����t-N���מ�k����MD��{�]	��F�<�W���d�r9�{>�fjr&~���R��OC�Lr�[t-Oi���/0G������0 ��P��{�h,x�D�{� ����Q�����p3S�/"3�r k��L��z�B��.�Uu��;����8�G�:��y�-ȍY;��:���{N���� s�ݯ�=$�;쳄aGĄA�K$�&��M��Cv�B�-?jJ���I#�׏�<j�����n�<T���mq��2XL��.���e�-H�CږQ�ZֶV��庀�������AS�ˋ���2ôrW=>@��π%<��a7׿�}�X�T��t�	�<7m@}�t],�so�,�z��Z��=s�~Ė%�yFwU��i�~~KK᫿�F��pq''m�M'���aF�y �>����xla8����a�ՇNtݬ�?�y�)l��9U��q8�4M�n(���Oj�����2{��Y|��ޤs$Nᛒ�M�bd�]TW:b;	�Hm-��"�F���TCЮ(�}Zh�w��Ҧ�� \����}�i`g2�����{���c.l�Շ,V���*6r�����:��x=��������K�R|������\ˏ��t�:ĩ���݇T�m�;���2�3h'഍Ml_
���{���(ˆN�k�+�R�[��k��g+ Z��{���v4��w=�_v5�mۅ�lNp�GG�)��t��vwo�Ą�V9���R�.�؎�������^�#fe�^���"�m���ɪ�Ƕ����Y.��0"�7�k�67��v���a҈�`�Ϲ)uiD	(�2)T��m[��V��?	a�T���� a/��c1���ރl���!���-�14�Op����%�4r1�b2$" ��#Ð�=틝�N������8P�̋���!�I��:Z�S������kU���D�Zz���� ������58��J����'N둫IYʟR���uG�>4�ͦ k��@��{pe��:"\?���J�3`�cG
p|�Kc�s�6�ъv��P�Q����)�h�����l�o?c|Y�jv�l��;LC�ir��Q��8��'�L0	?
H�����0SW���2��%�E��6Y���šd�W+7M�r9b��_�����H:}GOf��NI?B�ٯ��G^���Y�O�Ҷo���X��:4�UF�������}uP\��� �@��,���\�!h�����Hp� �]w�g� ���m���}���������UM��{�O�>�9�ӷk���,�����M�b��Ӹ������d�S��6ki�k��lVh[���D�t���Nbp����2o���| q+��=���_�~�̌��Z�=�����e}�iY�E"�kh!q`tS����0��h�*:t&"a{޲pb:>�|�~˃�pM�0!%�y��5$�5V/����i�4r�^��3d���엡���̘���Svo���n��$�ѓ���l;���um��&��q`�|.b��lo��s�(� ���۸�*IF��2=�.�<w�㟃�Ҽeuop�i+��{5����>��PO}>Zp�.]�{����rhKYn��H~��_�l��yt�	(��'f��`Gr��2GԆ\@�}	�~�{ο�U��@ ��Fw����)�~�/�p���_ "�+w7�ћZn�:�E�iA��^F�5q3 �����B�ګ�E˨��Z���
^JL����|Q�n�3��0�-��I����h2n��*�#z��/�L�0&!9��u5��|��x��S����E�`jY��$s�%���L����j�=���G��9;?c��ײ��#����Q���1c�F7�;bHF�����b��	o9��T"/��!���q��P�������g�Z,Cͺ�f�°���b�Yp\a{��/Y��CW-���Z�]=��#`2�rA��/���it�@�Cn},��)��b���ݳYϵ��K�/��V�Q�*�E7�����w"��bx!U���Y�k���|���W�]"�u�T+n���d�'3�`#��#��<Y5&���@�a�V������(�u���9ϾI}@�0V��{v�r!�<u��
�X�	�����tB�jf�@sFqsg�rm�\�6��3Hq6��0��zs�}s=�6��v��%������z|w�4O�a��#�%u����tP�������ї(1�w�޲�i<UWW�t�"}��5��`2����}�T���|M�yH�_B^�/��G�"L�\��钂��E��@U�8�6�쬝1�������2��1��R�d��=;C�fn�FEo�0žMf>��>�0�����ȶ�]��'[���?�ݏ��=to�� y�����Ǆ�݋��$����+��\��@.�Q}b��Sq.�t����  �	,��� R=��!���1W	8��B=(ȗ����Cw�MSz��TW-r�B̰������F�Q�mV���{�c/���b�.ǹ�7?�A�
�w_�<6k-�m��,��:CdF%XߎN���t���qzɒ�4x�q�~�]s�"\>�QH |"�<ڐ-j�y�f �����"Tט��d�%�\��m�j�ؿ�� ��ku�f:�i��>�!۱�rQ��|#��z�����(���3I�<�[�,h�*#��F!�<c>����
㥒��xw.Y=�zFҝ���]� ��;���� �`����&Q����ql�v;B/�H	}�]�}�ؽ�! ��S++C��[y��H����D�����R��k��M#���)�,K���7p��F}Su����}ڭ����K�CPF)o��e��'��B>:�Vs��umXg̍�{֐(�<QW��L�^Q:����o�AD1��L~�.���FF=���yYc����W¡�����~��Q�}��b?��gR`/�H{@�1�K����O/zh���������8�Q�5,��$w��B\�и����M�+dG�7�ӯ���f\	x[�mc�$F����2^���T����q��0|m���I�^�l{��C��r�ƅ<vcᅂ��R����گ������]K�kd�}�kX�U5�tq� _����w��@c<]���+|�
��;zF���e�[���d$\!H<���)���a�W�q&!G5����G�n�0P�c}����_
	��z���4xЮm�ȜZϔ �u���4��z�"���(���H�o����,뷯3>�1"v�}��An	�O�??�l@%���-�^̬Q&5}��֏JF�<��,���ݍ�>�ag��ݩ�hi���
�=۵ȗ)�3�L9�l��9��g3�JfS-hS���i"��D��w_���F+���|���5*����F��/����m��Lu����9��#�Z;_!���I��W@��;���ɇ�.�ծ�\n	ڿ�:^Q�u$�H�lxLr�u(�����e���ϼk[�$���s	�M�'��TtOh�u���]�k*����#'���]�P��0e�1
�l��ǹ-�t͎���h�����ϓ�ׂ����"��<���@�����6&%a_[+�8V�ݸ;��yr�����϶|a��k�m$��F%#8�6II釓X���S�=e��7�L���O�'O:x�
Z�s��o"�<x���Pd�0�������67&�m����a.J���%Yc����XH�k�.[*�H�y�P��[ِ9��!�n�	�3�Q��^��G\�� ���!?D���"��1FQ��5�>��,���E'U�oױ�	G�HjJ�צ�d�(�"I�K�|�L#� &�4�#�F!� ��S��1�~4��h�P�Y�o����ŋ��T]E<�j���� !��������{�9�гLK"�:II!RW�iڌ�ց���)���}����Y(5Jܮ��;)E��؛�7j��ɻcAV�qH���Q<;���ݲ0�T���܊tI�s:�5��c
R���֋[;����4Oa�ň��43� ����ත�ӏ��ۼ�����,OXD� _�Z>�f��$�T�SX�h�|�;#sn��#�]Ё�ΏB��9��$�9��^�H���'��Jί�\_q�� ��h����\|Dy�F8|�@��n�3:�Z�A֋q�N�G�!�|�����PSt��5c�XYʐ�c\r�6�����7T�Ok�,��R^�'2x�O0U���v�1�Oy5�o��P���tLb2T����\L��6Az�����"��?X.�!���E�2^[DL�K���§A|�'k�f�:���\/�
�m�P����ڽ_$<�*��}�&]y��td��A�h�f�c�˚-��z�D-:5D�u-s�pa��߳��HO:9'��j��~\Z\1����M`f"������ZD�اT� �6#~���I��9� �s�+E���ƽ����N/�s�d��y!��,�R��8�$��-I���h�埿Ĝv�%��s|G"۬ �nt�c�ap�)��-���O�A��è��Ǹ�'����lR.cFو#����]�#��l������*G��������bO|�9����鱲ӿΜ��[�pb�=�l0+�q�R��MyU̵��A�,a�og��,����Ј8j����j
�^R�o��uq%���\��tWLM!M��sV�ar!0S�\�������HH>�Zl��e����=���Y�ǘjB��I�c�螣�l������>3�C��a~��tP&����|�U�ĸ�"����j�6$�x���~��7b_v����C;ơl9vC+��Ga|�����a�����n�0����ކ�X��yD���h�����g�Z�b�Oq0k�F�z�U	�n�U�k� "
�!]��v������ټp{�ď���"l���rr��L�� \\[#����;x�� �%k�1 ;"�>�O�|�'h��|�刻�5���o�}v"�,�RB��j��� )_;3��ʆ�eC��6eN�|�I�^�m�~� @�>����Z0���L	)b�}��=�×���TR^��7 )�d�ѼP=�l>,dˏ<�?��W?�$�>�7���?����Bn� ����,�z���Z���u�H\=U<�߇���c?��uܸ�?&k.m>�����_�$��@���R��O��� �eT6e bTU����2Q[1�M��y��ӷK>�� �Ԍ�i��I|R��c.TC���__�*��X�yX��9�&9��!6���-��l��s����rd��7�Wc玠�qe)#��7k���t���o\��l�Е�3�&xV�_s��u�%;&GI�.�@���c��}���EZ.���.����
�<�ā��5���!�ySн�peI� ���D�Y�:ą��� |*$�3�e8s�4���l�ț�K�Y6�@�7$�^6�I�$s(�	>@��}��0�4Vٺ�|�o���� �{����$�l.sj|*FbN�a�HaPm���Џ(��3t|t�"���,1�ow�MRN�*�0Q�Iu)�;dl[�J'�'�k�k607sw��<`�t�K/%���+�E}�������[J��� �B�ͫ��ӿ��߂Y�O������3���prLXs4�X��Q�����5VB #�䤖@x�{r���)�r(����am��W��F�\&�$�����]W��ݿ����D�$z+��������uƯF�ۮ�K�(����^�{s�l��Ǩ��u,;�ˉ�j���]�@-|�^����=l�9���v"�,Sl��C�����D����� ����Qkҳ�`�ʏ�,F�~�����FA\�VK'�3�ԼK���%P��A�A�l¦=�jf�g)*v�{�#������QU�
8�w��c��a���{V�%P��(�Qe��$uU��d���R�����|�����. ��x�X�' y���k�Hցtp��ˌ�'����p�|̵��#����<Z������˰d����}䠌�8V3n�!H���hGM�2���27�#h��#V���on�a,h��jx�>�\\��9G���3�r�԰z�� ��=�_�����K�ӹ�t�N�=Q#���;�?ta��_s�����T�+L�8~?U�4N�1�f�H-x3��H�����G��B���i��b�/��P�r�"O�IOUI�`�-�S�Dv:	O�^=~4���?mp5�������G��BA]D��3������4FY���$"W<�l֖�TQڬ���~�m��<�W�uԫܵ�9ֲ.����\�$ys�a.&�d�h}{v�w?Z�s���:ь���7��)t�wٌOɱ�myɢ v?x�t���O0��*��_���cި�l��x!ٛE�%�4d{�y«����u�(ZT!�W	A�^Ѫ�[��;�?Y��kj"�#��7Ğ�އ�:���1��o�j���������%V��}��Ml
���<�㌕���2.�J�M1?Vo9'�a����C�j����)^5��5�D?�F"G�c	Se�F��t��*6�[�Y�7�>�/锨GzN��%�!�Q�lB,��VYz��Z�V\�ŭ��O=F�>%ƣN��o0n|^������u��s����G]�����2u_2��Ͻ��J��A�\3slydX[�Z�B��<<�5�~v%VQ]��%�:�+�e��|�T�:<GLC<AT$�'rzП�h�M�̧[f�e3����DO������
(8��v��TWy��k7̓JҲB�ݡ�D@�C�V�]��X�p����|�M��$�/�u7���9��J��M�~KWm���H*�z��e��2���2Y� ����� �~�Y��vj�R	$�ur�3��_�J��~���<:� �G��c�40�j����4X�c��y����z^�!�Y�1I����ɱ�HQO_��j�����bm��i��$�Qܘ,h��l�c�ss�s�d7n\}�)$�z�!���k_4YL�f�����h�g�
~[�F}���H��� %�<��§ˇ9�	����e��͞[��t��3�'���J��N�'�\!�l�����J��1�{.{�Ѕ�tbL�;��b��?$V>a����=�<a+�:�|p#���(s���X,�e#��x��LIs�ni�b�����F�'�����G,<��1�R�'cZɕH�u祪����q|�h���c8=������`Uc#qt�v,R@t�dj̾�ygb�Bp��:�N4�kjCW&k�b�l且����,.E��o�{,\]J ���})OZ���j�`ZS]
;�����˘ve�l����8�#���
Mnd]WUGbm�qe9�4s�]�H~�>:�:Xs���|,)l#;m'���p�g�����V9Ä6;I�d*�r�}�CL��No����_ʵ�bt�@g�b=b��lNn�!�S>r���]�C�5|�-� ��6���e>R6�m���t����І�S*��lG�J������9���w+�h���-4�jYQ��r6��Ao�������81|z9v���[U����f��yW-[W�uu�'��=��������6�� m��-ɀ T����J/V�W8��P^-��H*Ӄv��=�Pwf�{Q���F��X#�S��Xs�����F�U>��Q���|�Y��g�H�#R+�^��+Ħv�H|�]���+D��.��4mY�t� i7�(m��_}�jia
v>#]`��EJ\h���c&�կ���Ӌ��ST��Q緟����޻1�Q�C�er��-�io�@�����^�k�Rʧ�	�:t]�'pz �t\��Ќ�X��Am�P@��4v-{��:J���r��1%/J�UF�薌�U�T�0>�����8����GLu�h˨��k8��q{	^�͓6djr�I���_�=�Lx�p���i�7��F�Iv��b,ݾ�����H��ԕr�4s��X��V�����6/1)X���5a�ALӚ��n�HX��D�9v�b����}`�hf|���6�Pb��Sί��#�IR����7���^T�Za-d'�7ޔ�D�Pr1c��5�>Z��4h�HciҊ���:!NV7�n���bT)�0����.���	���P�pٗ�^
!ڃ��}�_oȝ_��j��qmӗ��� �J�:S\6e���n���j.d-~�'8�D�{�כ�IϪ2J��h�M!�C�.��t�;a�,������R�aHY�����	:��5�y���;��))�D7�\�8��/n��c�)L��z'����©(�W����c�g(gn"�J�&ڶ]ZFO����${�_E���\	cz}��v�p����u^�7 ҺA�"�_�B���*΍�t=��؈��H��U�%^��������a؍�kT�a#F�e5�-�U��Ϝ�� �����pz���6]T}�;�M3&�R��8�r��ю^�",� ����J+�1���4,��ňȝ���}�g�(%C�-N��^����Qҧ��Z�X=��Q���2|M�.�'�d��Ӻ�6��T��И��3kJqqh�J9�� B9�ƛ�]�F� x0k�)����z�5ZG��@��������%�F(ӟ���괊b�#ڬ6�"d.e��w_�Ҡ�-��_�d��}��� ��>i&�Q����8�V�F���d��_3	����vA���&���ۆ�wD�&��_�˸l˽�px�$��U� �d��d�"��3��u���D��j�"���[��˟�y�rE���(�6�	J��{&=��1F��q�V��c�DůT۫��st���4I��Ih�ؘ���LT����C4e1�gN l����,� J|������� �&_�Do=�,�0B�j}�VƝ,�`y�����X��[�ݩ��Q4�$��=�9�S��%����;`��6��y���4��܎k㥛q�+���D���������wH/�����FZ2u�\�8�(��+�<a���>��wkz�]�|�24�P2��ɴS~�n��{{
��J!,�|��-��"}���>���pA�nS�q���?�B.���;����?�Ѱpr$��L����*Fi���ѵ&51$�	pY�ܵ԰�I1��e�5�5�meƖE�	��U��̯j�`��v\>��ʡ��%-�y�����ohl*I��~���񮙴>�Iw�z�@�jO���y��6Ќ����h��L^���un�YkO�;�u\�z���/)�.����v��	��&�v >�^2��ܫ��
�ۚ��y`z��3��ZJ��`ع�p�lC��7[���4OY�lC���|Z�Y���̴��n��?Rvm<|�M��:�x3n��V�E�|C�g�zK;��r�<��wB����y����LԒ楱�D�˿�T)]K|ܶpma��}�U�Wf��350�0��~.Fu����^�Zg��[z�R���T|���l�~�P��%k��:֟�`$:<��JU_5��qP���!g^^�d]�^ټ7PH�6u�E�=�"��{=�	�9�<�+���:��u\�pr�Yw\
s��*+}�8zd�Au8���w�圳V��Qr�}���	�裣�@����vt���jۜM�����j���i��~�2�<��S�^6����;�m�1�X��|��L� my�a�2>n٫` �~����Ί�-*������
�l�a (S}�Bo�R��k�xN�k�h�m���-.��LK���S4�-��Ĉ�'����>q_WY�~�ǑC�c��3O�����u:N�� ��,�B�'��G�ۄY��fޕ�b��I����M�p�����N�����F7�����n9�mY���
�g4%59��T�# ���¨/_l�[f)/�?rEm#+�Ve]G����we��IFyP�Q$� ����p>���ŸP��X�F�����h[��ca�M�
�tٚ���J���D�? /θ�+� XW�2�l�o�:�A���*��m/㗦:[����HEEE}�����I]@��򍍩eZ��L��݌]VD���>0���!�������d�SA���3?V ���f�к8k�(�z� 4�� ��Mc؛��!f^i��큓�d�tn}T��Ҍc�<\����:�0-�D��H:�\�%柹=P%%�9�n�F�YZ�(�F��Z�ݷ^d﵄5x(ʂ����G[�9�ֿ�,���{����n�m��,�j!Ro��W �������X��3cKxy��(���=����L��Mɤ�w�x�?�!�@�Ρ(��m�T�^eL"�]d�G��6�xI!���8Ջ���>�����{��r�, <��@myi�Y:@	
����y"�ܯ�~���E��=�����y�غ+le���|��1�?VZj=N�lڕ�J�v�T��9�_6}_č����e�9��HlۯS����g��{���Fa;At��;�r�+�{K�QtG��H��v,��D�P��{�O{�Z��%�ޔ�9-��"o!3������\���	󖥽i���Ӌ��xN"u��}x/�$�2�<�2�D3�u�''����!�k�V�X�V�WB �*nup�\W�����89-�N�"ô����nZRE�I����}4e�*���;R�"��-x�[��Alm@l���OGL/v�5}�H��K��XY��Q��s[W�¼�����ڒ���ӳx��Ṥ�M0�(y��j���}�´G ��W��k�J1{�)���{�`]��E�ā�_I�m�ź4�@��p<��ɓZ���ɕ������`,�<�d �"Z�)����E6v%�rޜ�L�\�} Q���]!0ͱ�B+��2-��X��1���u���"��6Z�($�T�;����t�߭|_�N����i$�3��O�zRƙ�@"J�ħ~�h=�g3h��0�Q%NZ�Y~���<����E���WEo���a��`����IZ�>��m��dQa��EF_�[ L\�{���5���X��-Z剁cf��L�B2�y��S����we*��޺��9\\�A3�z���P�Q��6=�͗�ע99a6�2�K�<�̿��4Íci]��x?4;{$'�g�2���������4r�en�m�]3��8����Ȱ�j�x:.�L:y��	\�4���)@��±��p���v>�ϙm�Y�%5� S�i��]=e��-�*V@����!�{Q=*�_��5�mґ����P9:.Ňپl�q�>�Rp�8�t<�y�	M6vNh�G�~4�4Q+J����a���;�6w�_+�W������;2uM�\(�q���D�w���p,_ķ��f�ג��Q(֔uϚ���3�>��x��	�R@�����.�i��զ����W(ߧ�E�\V)0A�׳�r%yP�1 W�D֘�Tg.�L_O3i��R�~%����æ��mڤ���T�˚�}� ��ѠOPv���Oo-�0�"��g��JWy���r)S'M��fO�Mx):m�?��*�ӳ��L�Q��j��M�~�H����Z�1�."@�����OZc�z�:ur%�@�HՉV����K�����3��)���X�_VˋN�JE�\/���w��1�_���eM<�箵Do�
}��_���M�>+L�t(��}��'�ʨ,!�\5�N��ĥl�閻�]
3*���4p�� ?�����i��F$��%�J���A�)-��x!2x��vt�r�V]]*BS��� {5���{`>���[�����AɌ�I:+ډ���D,�6q��bx� U����l�+�Lx]1�F^ţL�&�Z*UF�H:��&�<J�H<�ݨr� ��T��nCݯ��+Z�m���<
"�	ۖߧ�� �<��樚w�V<�gʸg�~lc���n�=AZ�PX�ݩ��VIR� C�\.^��뼤H��D-G��o���
�PNϪ��
�@JW&K_ֿR�/����3[��׋TЋ����S�;G�ğ��&_Ud�Wゾ� z��n���=�G���x���ޏ�t4�n��

�[Kx�#�H���) ~����{m�!����nr�dv`�9�S�«fL�
�k3��o�G�qt�u	˴J�j ��9[B�.q=~W��S��T�T�TӇO{Ғ��B�b�/22R:	E����I���41ɫ9bP��q�����|m���0T�����G��a�ܪ��	�Co��`����:�2��v��/767M�ޡ���� c�-<@T@�D]]]:	���fO.������t�@0J���3�q�ۅz�5� ���LQ�4{T<���mc�g�WyJ��8������4c'�CH bO2s4���f7���XȗG�<�����][�;��	
�? f�3�OK��/�a��/�QJ{{{�=���ƈ�qNzM��_�TcJFFYTT�̟�=PƷ\#YQ@����]��v�>����&&&�T���dW;�oQ�uG���%I��)�l��< 1��͂@�0UTD�߆NO]�GFz��B)\���,�B�%2nb��XP�Yv�`F�D��q*AQ;[�R����UH�t��X6_�Л���NwB1�@+�0w1��&Ahꙛ1����Q��)����)c�v�ˮCA����v`&�W6�܉�$�)'^�����ܒ�T:	��4933���j���T+��xw�i7��I4UK����Rݨ^�/Ta�%Yg��>�뀥��Ol�:�$@�VԎ��/���)��Z)��Ajũs�[-ٔ�>���]���~Rյ�Q�{�Yiq���.���,�$�	9Sn��"�=�a"�B� �џ��M
cs��3�a�������Ϊ�vِ���f�?e����A�W7�l��ˍ�$��ocs�,�5����V�jz6ɰ�%ft�#�B�9��	0����4������l=W���ͅ�X�	f �8���t�?b�.d6]��߽w#۩�sz!Pi��,U}�(�����>[�# 9��=��F�L��fd}��F�}�!F�g����Y���5�[��}?�
��=\��չ D	��̳4�ET������G�'��G���&�:8r�����%��5�;��
�Hf�����c'nTi�Ǎ�����=}Km�g���4���!+�a�m�,����������ڝ�݊�.R�.l�p���}PwQ�6]�Z(sR��t�o^������B�]�h��-�G�Ӿ��ck�nުT4�8��f8���)���V5��э��3�	+�'v> �&8���?F�Ds`3D&W����eZ�>b����6+��<��ِ�|�Ʌܘ�f
�LY#q�u	/���c������m��&''��<�}lDs��IA�/dc)Y�o]�D�[�o6�����ON6)�oL�EnVӮ�0HҦj�}��#6�����-6q���#� �����PzU�$w](={ǣS�ot�¿��06c*�a�2�G�Ϸ�(����J����P���3�ﯤ�@ Y�M[�h�.�B���ƀVk>��0JdF߃A�x �ݹ��E]W�o�F3�0���⌇j�әCJ(�ܟ �0�j�'�Bp<bG�k�U�H���c2*�Xs�W�Nx�}�x:�*Xޜ�I'u�����P=�����AҲ�@+���#W-Eq*�$#?00	Qa��y~oǓ.�'p��P�X@�L��Uy%Lፇ.h��>���[��U�o�'5��B�bb�fgu�f�+���88L����۱-p�z�!���E�(���X75�' �C}�#��
8:�/J#��H�@��)kNN5�"��6�ss��^�|�H�x��|�U�#��Pt�i(��p����e���,�u���	%h�
���^���;?��	�� .�\F�"�B$�� *�;�M������l�ȯ�Xf�U�H?�q����G_���3��M�~�)�퍒�2�2=u6��Cc�*���)�h�b�a漠q1{|\�$W+zn�&)��x�y��Z�$#+�9�ǔ5"V$�yqwP!�~rԎ�d�?\��w����Y��>�����	w��~x'���M�j��wL����Ӏ��P~l�p3��)��눿} I��c����P�Sh��޿���6`%0O"`� Ǎ@�,Ć�p�p u��Sex��P�
��>���g�$�4���yT��Օ�O�����Fr�d(_�t���\�ȕ��+J����Ų���Ñ���{�ր��_�t�����-��Xހ�b�:|/`*��o�������n��'�N�
�c�����Z�;����Z�8zy�'���B�`i�G�$�i �ph�?�x{��G[8��H ��Z��ؖL���aYtD���P����A�}�{���p|����b ���|��<4����t�x�ѽ��{+�	�<L5��!�W�}Cd���b:�p1೹k���g�X� �{\B��]%t�2�'\���>���:�'�B���}/ ?����`�p=�H1�N9��h��܆Z/�J�/Jh�����V�؀nm����Ø�w�ޥ���8������@�q<{�����!"b L3�4$@�;skn�Zl��UYU�9��Ks@Δ��jrA�"�նv������Í�Z���j�,A����QM�U���<V���}S'-������r��:���:�|FnO���B�Ր���~cw(����	�E�D_0�\p5IUӗ�HĪ#�iGu�,�ˆ�˗}|����T��gݟp@����K����*�j��k�ɮkb�G�Շf\�ԗ������G��||f�'k
�[ g�y倮"+��Jv76F��J��8�e��T!cqqq9]���7����9mfx����iE��%%��/��������Z�e��x��{���$����mEꅫ.Y7��1W�I-t�{���i��<�[0��~MCs�p�C%f�(}���Pΰ�(5���D�RR�c�5=�ש�ot:� �3�^g� �w�[7��N���tP����\ŀ�����F�q��˓x�T.����@dxX
�0Yt_st���j[�$\\�~��lu�H�ca��嚚��_�,�ѽ� �T�A�S�҄NN�ņh_A��.��Q���%��NΞ�y����X\�-W�rJ�&\�F����;��A�!�Z�w���FzU�Ѷ�oZE���NW<8�h�5���@�Q5��.Od�ӳ�o��|���x�r#�fLƌ� v�V����:�����&���ɻ��N�z�������_-Z5@���b'��-'���/)`J�/���D����^$α�}�ȪZ��__igL=3��f�c��(�����v�D�0��ҁu��}���rƑ��[X�`*�;ġ�6�X��k���r���*�V}t���^t|V�3777p"0��V�c�Q�k'��)��:g;h>`za�����ǔp?>�� �hih��=�ճ����'�.�a)�L�F����	���4�ޕi�����~pu���'(6��]E0qP�qB�3���hc�4^'���-d۷4�h��ɺٹ<^�k�yn)��VQn-�]���yk�x,�dc��<��"$"�&�xK�x)�e���/�1cb#
�Ca7s���A` c"����uY(����,�4i�*�뭸�x�ƌRE�9,���
��WЉ���t������]<u�|7c�lA��w:�����Ɩb��W��L������׈����B�g/�!�Ev~�t�������s�m.Cn�]�p�ͺ �}S��Z���ϸhl4��q�nD�����U�9��f����B�.xd5
�S-S5�9z/�_�7��3�#NV�!�����GB�T����������kGNg�%y���u1���K�BM|�N�\m;c��G�ط���.w��
�\�;��d��y�;*�Ǒ�)4���ƾ�^%��e�uN������?�,1�#��k~e?�޲��"2,�k\~/E��
W?݈	�f�����i:ק6m����c������͢oV��M_֙Y���Ӊ&�ş��:z@��.�6�z^a�'��gzl�|���Uԫ+��h�<&�d�w�-ܼ-��va�<@9⻹)zZ�����C�EޢY͛��Qw-�Y�HwL�mx7�ל�iY��Hh��ն1. `k:�?��1�k߽�i��ۺG�LR�ݵ���i�zb�s[�O�tzt��&V@TɊB:����j���l�{W�&�$l��2-�K�ܧ��4<^ԁ3�����X:I��1Z���
J'����}m�t����"rf��zV���k�Ǣ�k�wS$O n�;��������'@ٮ���.�J	���my���j����e����P�5�*Q���hV���(�d,����`no�&´/~^�>|�o���"�:�`�~ӲRM�c��|�u�Sf����t(��h�ݐ*�ȫ����a����!�q�!v���s����n��r����o
!t��H�@��9I����~��aM�<NK���y���o�h_1�����	�f:����
j���=��w�G�T^ڻ�˺��d]W_7��c.C��C/�;~��r�O@ӈ߃\^�%aj�,`�2���i+�;�~W,d�����[u9�ժ��L�!Jw�EԦ��&z��{&T��LN�*�z��uW�
��/!{������<Nl�cp�|_ޜw���f�u8�����w��>H��W�Q�%�oc��-�n��b�Zh��ڭkkm�ѲBq>�GS>�	�_~�/ �ݥ��	~�,wqq���B ��Ę�O�~���T�6+�Z��*��w����gK�(����(��!-�.�)���D�|5�)@�3�]Z��!�Ͷ�]����8�_�N�/8���'T�������M%t�j.�x�K ��.�g׶�l,e�G�j�`���yD��Q޴���;����}�]�(�ܙ�n������\:*))I5sE'37s87Y/h�����<e�V�o;�;�2"������B���V>U*��>�	 �mG�RR=(��8��
�V^ˍd��)ozIy����̘�u�y=v�x�Yc2�R�9�4�� ���}�Zg8:�5*�N%PI� �\P��M���Œ����'�(���"m#_7}�����7+�z������������y���*b�W�n�xNK�ET�_�m�{��VT�U�!1j$�U�?�϶����1�7K�X;͙%��%"vp�bc��f���v��[NF/�g�)�c�8��ʭ�{��!;.�b�V�}�"ވ��T�H�ڴ��l722�h���Qk1�Gh�#E���ʘE���_�,~#umQի{����Ô�D�zBH$�`է�1�ᴲ1=�')r�t�-�e��P�*@�̶�z�zX��5��x,:�.�v��S���<:u9=�;��;�{W1����xd]չl����jg��F({�;>,r~���ț���H��H�̴L4c�^ Wӑth�R>�S�Hz8H�1�6���cQ>Ţ�P�;�����d���h�r�)���suuu`�k@Kp	���RŢS�����lo3��(�'T�Ƶ���{�|o> ��My1���:����'#UV��$$�^�~�R%S�d�H)J�Ȉ�����:���=�n9���WְH�F����VN��!v|��,�� ��7=L���5uĜ�4��V	Ԗ��Ą����g�V���t�zw��'��~]j��_�-#����|(�(G.�'.GBF�@x��YH� 8��  �a���v����o�O�S�{Dw��~L=�@�:A�f@y��B_ӌ�ׄ�"��|ˊ����ί�c`v�e�����~���e�:�ug�b��}�v��@���H�A5x�H�O�������ɴ �p5Ɯ�}_k����D���(�`ut@�w�g|9Y3�k�۪l�����Dћl~�e�iS�U�x;�l�	 ���2�>Ûp�s*a�6�� /�<���N� �@"w����X��s̒��+�%��_���Wqe)|��Q��
��F�"1� Q�v`�vW�;��"�0�!�}c�h�C�k��=uY��"l��w��]�n�h�d��k,>����P�b��'��:*ʮ}DQ��0H��nP�i���TI��n�T$j�a�����w_����?�Z�Z���ϵX׵�}�3�c�=�.�5��vTA�YE�w�'>�oK<@L��ۻ2<p*�k������#i��>��@��p>��a�e����)-��-�hs�e�NFUǉ�J/>Jb�X�����m� ���矯O��L�6��R�l�
s2�zc
S2���~,�~�w�N�=8��1>L<��i#�fF�Gs����7���f��}��g��=|�QUQ-#Z!�P����E��{&�������N�G
	?1���H�@�5�,��ZQ����Ѡ���(�:SC�k��j$�\�����9��)�[�<� ����� ,������#��[v����d�k���`-�;Z�?�N��c�V��mb-)�����o�|�(4�(&O�?Q����s�[�6Fg��Vr�[��C/�aZ�smۯ���HWM��s�7��������N��9R��])����`����ɋx�ߍs2 v�A}�#��ۥiq�JGD�c���{�$�3ְ,�����㝬�[�� �H���x����e�c���0�v���q�����Ց��4���|(;���`
�$����ߋ(�0�Xƙ�85-E� tb'>*����?�֩&��n�Q�	I�k%tLG���+1�B1��qDQ�1��	��`�b��A�5 �@��q�뙋2�Up�o�g�4�V,��	�zw�}�%�}�l�lxs�M��kn �Pl�o���Ұ�7����ۙ�_r��;h�~
bD����. �XI�.$�B���iՄg"e�I��H��T5.�.]9D��e蠸 �,ji^�U*2�=�|-G#A�o��S��<Ya�����҄���N�{"S+��@�R��b�2��-c0��ޞ�;\M�W�lL�+ְ����v4/s�3&UѸ��W���9��UN��FMs@��/�4���ݦ:@ݚ��@�ħm�������6gE�@6�����������IA>&�>���kaʎ3{�-xBC��<$��qf� m����T�-C�۲C������|��^50�v�hA����_����-Ƭ���Mm�&���xF�ã�o-���&\�ui��~�_+_ 2����cH�C��ޏ��Eui�q�*�}J�H`��Y�5fB�x�i�A�k+@��"z5��2��
U���)�z�/���P��*�@O���(��vf����+hˬs~������NBbv/k��}9��I-�:�Q�� b��&�G�-uZVM��	�������4S��	(�!�l4Sϵ[�m�I=�S�����?��
�U�6�[|�˔���^A_K�Zoi��i�^��xkN:�Fb���7	j�a�R��*<^�*S͋�/�:�0����X����vȎ�i�R��#���ipL�y���O��&@��W�Leqׂ+D��ZMXO��4�>�����j�tdq���eDߺ��4���ʖ�7*WNʳ��S��>^���G,��������3>�(�wF�l�b����1�,�$L��ȟ �L�`mW����]���i�9�!vT�,@��d���ŢM��"��Q���Z$�q��|��W>^.�(K��Z��?Eh�h��K݃<4�Q�^��0�:b!A����N&��M�f='3�wV�qhh虘�C4^��
,/�gE�tu#߄�_�`V���%Y�c_��SϮ�h��="��퉻*~u�E?��#{d֌Ú��?�tb{��K[CօxA�9�"���)Ez!�"������_��D���A�J]������Ev��-t���w��iH�\ӧ�^���v���{X7W�ρ�\�:�;�����pvj��o�x��8�=~_�Qm�&�����l�O�9�t�s�˪�ۗ�%�kD/����0�� 콯�z���M-��{�\�kV_k�FG�Ц����8^����uA��Y���77��m~Ԋ����a�/��0�H�&���7�<)�ìYv�
�d�밡VVK�u�;�u:M�wxdj�V�	�ȵ��u��0~*�~�q{�V��ap�W?��AB��T!�/N���R������������ϴ�Q����)�4\J�ABS'��?[W����g�ҋ�x��k/�'&������k��ξέӋ�I��NO'�Q�/�<3v
r��c�w�K.a�~�"������$�|J��DR[Sc�u
��m{-z��׮2�� U��C)�W\�o��~�	�ě|.�8{��Y��֯���fhΰ�f��$"uq	��]�#G���˓�e��gr>���v8�z����!��%�{��mu?��W��<L���Ƭ=�/*�䫪[mJRI��Oe?�l��٘1��]�C&-������a^'c(i)�,ef	�Q���:<�-r~��yZ�~���H�T(��s�C��I�#`�Z�`�@�ܭ��偁��{���w��۽�p0�L�#V�&��RƘj��3�1M��݆Me ��>�;)ٵ�:p��CN��϶�D��eO��\�^ �5�;	#;O�6gLcD��p�y�[��'�m�.�������^�!��������{cʴ��%�߇��|����r~��[���b��;y����#ޮ7�o�i��N0�$�\�3�����kQ~^���F+�:��f���S�cP��Eb�,v��Q$C����$ʞ�+�3�fo����[+�����.�(�A�I&�Ȓ��uj��QSC�DӴ�B��$�q0��-�'�,��~�&���T���rg�_�H�(���B��"sv4�0���y��_����Ӗ�ym�Y�
�Sf�SK���.����^V��'�+��viniF\8��-	;�Y������qEb�^&`�[po��K�^?;*x���5���߸������ k�k
�+/s��k���ՙ��'.�$w/1OA\��g��G�2Sw6�X����x�~c!�]�[u��mМ���?"�}�o�8�u-�t���#9����ǳ��/�<�����N��)�3�@�Ε@o��]��� �$�J����&o��X���<��Ua�	g������V&oc���g�N��y2Xn��T~��+�i�W]���(^1;_"��!V{�'8�"��ߔԒ�9x�k6o;/�L�M&��3�8�OEX�S�ӀI|�{����y4�I	���V��0<�r��F�u�j��q&����G���7�z=��!
@%`J>��	�&?��/�o(�U�Xv��4��U��FX�ȭgVS~���X������ړc� ����y���hqS��~խ4��?�c�]�����3�/19}��Tߥ�/�F�/��j�d�zθ6�sI��� �1J�p�"5G��Hɟ�|-�\��1i�t�Εs���?���Ա�1�̤�d����׾��:��b]�6���|���@th�j�|u����i�ω��2}�b����i5NhS'���G����Ľ�r�����y���iG���J�dyx��g;"�8oO�{�ߕڙ��cL�_~r;|�.^fֳoI4>�8��sJ��D�f��Ay˟Le��e�:7K����Svꙅ6����G��'sV'�8�I��'L碵'&��x岕��ʹ����/=���ѻ{�򘆛]�⁠Ԍނ����׿�.PS���,�ZMrJ�"I���ygq*e�t�Ξ�1�(�V�VK5��U��������Y�a	�`Ɨ�$`mV��2{#a�u����5�.+@�V~j���3�%�͜��S��?m��U*�	eƷ���৸���a�v������W������R��RO"Ak�C�}���[�5�s36�'�w<��	Y�_�#%.ua��$��Q�ы�o�!�̗nl���ߝh3��FGS��iXpǉ/�Z����tsv?�8k�;�+#Vj���:G���:YI�YؿIe���Q2bI�ӥ���B�v�uXO���E��������;,���nC��%;�JՅdA�T1�����	��pA��AhKa���P�������6���L�%�����%l��D�nڤ���T�X�,��,tx��x
��ܷZ�M���́��C�)�2�����B^�|�o��̀&�M��D���:m�����(��
����z��OCg����m	Y�KB�������Bw]P���MlRwSPV�T�}h����Ƃ���p� ����9�~O�_��mz�du�@���i����S�ى�K�f@����8�E݆>�r�Q�����+O��?�SRS5/���S䑩'��q)]L���k��{#O%���4�����X�c+�`XSrZv�B+԰��6�ia��'�6���V�+��Gz�	p�TZ�lAo	���mc�n���>�u��x��N�7N��	�凜�03?]���������c�Yv'� ���`�O��'��}ۧ�z7�D�<����`ƶr���NN.� �?��i��}�2X+0	ET�����i���d0�N��|�z>B�@�<+�� >ʅ�w\-�9�F�9.�B���Q����H'�h�
G�i�B�mG�Õ�L{J&Ŝ�}��a�Ё,���n����7�zյr}@���nY-�h���u�Z�<]s��_�ࣂ �ţ:������aۻ�u���m7�LU�ǝ�XG-�Е�NȽ��>�Uom�ή+�@��W,�z
-C	}�"O�'����؀	5R�gd���ni�m3����7�����w�7lE��(Z���;��"��j���"�C�Ⱥ&G �Y��T$�t�sU�cO����S�׀���w��jv�u�ݥ��\b���r5?7����b�����/3v@F���}�̸G? M��A%�d������̏-!���{/զ�/�`�Ґ�Mَ��D@r�Wȟ�b�w�C�p� �z��5���C �:Q7��젼U�N��6�4�J��į��z�~	�5�%W�	��J������y�Y�T��&�� �Оd'H������~Tq�h�0��/w�A�J���(�`!�?��6�(������X�A\���Ο	�?`���@�jޮ��=������?����y�D�R�<Jw�X{�4*�����^$��V�n�jb�W�#ޣq\#��[��]�:$��a��V7_�ox�1v״:�+�� �}w]ɾ%����XpA��w�ݔ ��y����i%`_ޮ>�T��g><�m`fB[��M:�2�U���c�L���B=3(�B`�7�o�]���44��d*����TW���ǏWu����mm�gΜ)��|8??��ãca�^��,����]Y��
C�a�Xp�9/�Q;����DL�3�� 
7�L�o_�\ �1.����Ұ�g�15����r�˗/�YXJ�ƞ�+(p��ܸq���J�ٹ�͛7�W��t������r��ƵϪ��PRRƤ��MM�c����7�t�0�iN\�l���n�qr�z^QQѺO�e�|���¢��$)>>5�.����e����.�=�r$h�*��Qe�[I����3����-��5"�ovޝid0�}�H{fB��
,�app�v�x���)*J���9�����x�)#p�,���힓���Ņ�B�Ar,�����Mv�{�	9��T��u�*���B6C�U]�򪫵�})�E%%-�;������;%��������|��r��U	
�6�g.�,����L?B�0;�g��|�9f��\�cq@�a���5c�&8���q��W��E�x.'�ZSK+69����W,2�S�1��Z�5�J�&�����jluV�f��.]ʌ�1,��k�'���㶗�>��_��cm5���2%�ѥ��%sYs�� ���B1*V\�8R蜃������%X/��ɕ�JfP����~=}y���4,�������R�Lpk��_��z,�Í�0y9[���������h�S³�o|h��rZ���q�ΈL��&B�?�DU�����ޝ>s�lQy���B�}��0�;u�z��[�q�F/=�g�b���4�%�Z��|�./\�z�W���DY���|��R�c�QWS�l�r���o�����W!��B�z���NSP�`:C?}��Bl&�����%�X���u��m3pw�[}�#l����5���v��w����S�-p�c2�G'[I�C(��/3SMI�<ΰۜ�������#�'�iov��#`��P��I����#��� �彤��W�6��/�?w{�%�^�c�ۥ�M� ۂ�D\�-���;������RTQ��(�X7�׳��P��R��5�ORFD�*z6b���+a��Ф�P�s����X���de;�:�<mU�����zUwm��s����)lYܫ-exDKY�W�B�/w��@2MW-��\����#��'�bO=,��s��]��㡦�]Rޤ��f�K��\������)�!�I0�q3X^���mĤX��n���2^Ƙ'��Rx���R�G��m������0��H�o�dJ��^�xE����p��_�$����R^n�X�>�b�x�qY�d���Zv���= <b@{��hV����
�
ڑ�n�r�-���ˇ/��]�?���z
6�LK�J���yR���=7e&�X����!�� �N���a �� .�2SE�����&�=�O�V�j�������m'��ˊH�~X@���L��S�^�u�MF<��\�+|wQ���1���K55o��*������J�N��r�/����
r,볥�;�� ���k7*:<C͹�D�k�e���X��D�d3�͊\":�;�j�>I�':��\ ��s ���9}T-�����j�So�{ ?qw^Pl^P��{f06�{i��٬n�c���9}��K�x =˥U��t)������'�y�,	����rѲMX�է��;HX��A	6�����?��Yu��}��²K�gk~�O�f�X2p�M�N�x�&"�� K��Z }����V��o��	EZ�^T�Y��QQ2V�xM��h��$�a�n�{e�S�q��0^ch�&�C�r�|��T�NZ!�}5c&����R���g�Gی�<�_��h�>c�H6;�\ݯ�'�U4�`��4h�2u��'�v@%�N幨\N�&�� �kU.��݂<oK�ͦ�E�p�=�6I� eK��M�暈ν�����1���Ujr{I6�v,��"�S�#�j��@\��s�tVs@��U9�b��ҋ�Lӈai��H�0�{w�*���{�Gc�:��V��7��p��ޣ�o��EJy���I�s	��}+��(�8��5PaQWZ�Q��&"_U���<<л��ޒ$:�oAc�2��G�1�dm�/<�?0�7��u0�U���ui5b
v��l�m�hg�[l�ppܗ�T�=I���k�m_2�t�`��	h�t+�wr4(򅼤��X7X�5��Co�/�׮_&zf0��<����KN*�H��BQ_~��-/a�����Q1o�Q~�\S�B���H�kψG��cvt
���݀�"y��6�G׫0m�q_Gm�~|����/A��@������Z������;����d��2���vX���3���g�Hi1��.`����}X�(�T�z�F��څpp}x�4ʲ�5�޽�JA�kj����4��
 F4.jX'�NIsNWN���߰aϦ� ǷYr ���%�fn����]IC֟��Pu�)�ef%��C3��A[&9�4{�I�? ��0����U�{����G�>�?$�[���m<��eAM&�����b4�4AH�d#��U��T}Bxi�����!/���m����0ɖ�@�ݦ]��xf���3"�]��������ǰ�	3@�w<��}�v~��3�c�y�[]S#3��鐌��#h���	_Sl�S
UVU�P�j�S��T�G�M3ߒ��V���|�R��v�m��Po�y��|a��8p�hWU6s�#3�`p�mI�� �T=+���V��^㩇��D�l�Ǐf�Y'A�2m%I��+�]Y��l�����eWK�(/Rk?�94�)//�����U*�1|�m�ܲ�?V��غT��`�rK�xtV�tOnas���Aq��naq�2�E��2-F>��F��G?��HP9�|�����-_�E��sG!��{྄j��z�͙��-���t�u��Wѭ��=�QC�tH\%�{ml�C�
G�tp�ϨΖ�'�ʸ��)n�+p+��]���`�y^Z���F?�߂{l�,x��H������� ��@˭]7��&�������$E�ׂ�r'����ge�G�l\n16kk��E�I۠,�7�$�� �T�<��	I�(�V'�,���B�̰����T��� �������ws#�]l#��?���zm#�bM;����/p,B���q���Y���'}�Ov�_��a�c���E,�M{��b6�Hw�>�,��T<�A��ON��BCߩ�ORwm�����=��$�:��x٦HO��]^1M�@�-2���$dW5����wkt�������&1?�>�%	� �~-䚥�)��%I�<�df;g#�n�xWj���Κe���O�_lh��ױ�K��6�W��6_f�/�{/3�z��Ӝ�mj���-�`Wy�.���PX[�2'|�u��ʟ���A^@K���j@����/���2U�MR8���b�S`H���	�*��d6�W\WC?c�J�����3g��8RV��M��}������}���x_�՜T�B�Wn�ъ�~O�y��Z�����&�+��5<��:������h¯H��7�}��o�7�i� &�E�� ��gsPE�I��i-����~�������QE}r��v2�:��Y��e|`�P���M��1��Zby��٪�ißV��|>G��l	אg���-�ɝ���Q���e[P�K��7f��:B ��T����f0��������z��m����׶�/���щ�)����ֽ����ۭ^u�"����/���4��жڰ&(^9��J���p��-'�98v���j�;~g�R�?����s����g�O��|s�J��ɮ*�N3�}�9�* q��9����B�-r��-���tr���c�g�:�t��%l��SGE����$���������8�hw�c�$�7�y�4F̭K����3�C�Q��l�������h�����<NM'�Q:�������?$�I�F���}c!k#}�s?Yw��~��3'z�`�0J�'�eOD��NA���ΰ������'2fnB�,�<�����l=��Շ�F=i%-�b�U��?��OV3#��?���[��ēW��<�ժ�J�_|nkR��6�%,u+o�������م�[������?B�G����'��<t�ڰ� ��OR�p��0w�S�d�4��>�/|2 �1�\3E��K:�I�/7m.�+C@����t����?b�|uw+ ��;|�V����7�`�&%0�\�dY���p�U����F�K�ýw
S%� �P}�Z�Z475�Rslk��( �H�(��x�˲J�@<'RsU�є髈�Χ?ے͞���c"��K�U��%��{�lYǛ��y��U�@����i}n_Zw1H߭X�&�KY�Ԑ��s�W$�>�Jڦ�}��T�c�+le�2��]�qU����}���K��>REB�G������Z�_X����+�l 0��3���	G�:������Tg�Ro`C���oV!��+ k��}���f���JZJ=�Z��z w��e�����1��mr�eƫ�A�Y�F}.�)ˢEY�Vl"���R��#���L�};��K���K�zm�Z�xtx<�x<=��� ;��u ڎ=H�I=�{�8�Do-�8������%�wrjt������{$�8��C�Z��-2=eBľ���������O	2`�T[�?�L���G�6�%�,^���X=����"IG4��M/����HF���7�9�y���t�
�.�5�ODW((TF&����>8x�;������DU���"@�$��c��߮%5��r�пv��P 9�'��?Ñf\W��lq�� �P�{�G8N�F�d���M�.�����cHA�Q�9�C�,s�5�M)n��d|�ғ��Ժ�CUd��c��֫�g<b���v�����uK�$�ZzW�}���;�	r�5K.[��D�/_������ݟ�=�@_�u�"�k�m�%�d=�˚�ЊOrwC&	e�|6���h����	�Z���]����˧��ޭ�p����e���9�TI��濞�[zI��+��YVK�&u#��C!�/��c��3�f��TN�,r��h$d��z��'Y�֮����K�;�;i:~�hT��S|��c���b���j��5?h�#���5��Z��qmv�8ȭ��{j����~�~�6�;�zt�0�8�.��b������`�]w]�;S(,���l;g��F��-�Lv֎��g���jHS�=[��8-�U��¢z�����Vtsy��� ����ρ;��TN�b���+�ti�}���nM�e�^T*ŉF��U�ʒJVm&���Ms���ԡ������񑞿{���Q�@�zԁ���$����N�{Ē��IemZC�����U�i�߽��yH�˖Q���On�=���=Bqw��6���_�E���_��-	0\�g����s�~�ZeY���i����i��U&��j��ޒG@��{I�yM�1��xw��f��_���k�`Wǁ(&/��H@6�9�$�����9Yz�)�aS^Rإ�tT�u���e A����#aPY���z��vu@'�v�Y]z	,9�U���`1/'���._y���t��U;��HV@,Z�X&&��6����Vb�^OwVY�Q�@���j����ة��r_��.��!��?[w��J:.>��[����1��	w,���(�Ue��
�"��y�ｙd��Pb��2���b����K�M�KA�9�%ȯ�Ye&��+
�>=�UNU-#}g�/ӻ��:��u6a�Z������^�����	��t֩�e����L	�CA��'}��w֚���5]%��O��"@�B+��7����VbV�VdT$���n�f�|�on�4�'ō�}�F����\A�βc����驓���� �BǿXtswB���S]�2T�	,6������@ɭ,d�������ĨeB)�;.�f2��.Z�5�����i���-p ��vF��U߳������E���`q/?�����)]ޒ��j�X����߹2��VǢ�
Z�$!x��j�WT�;��-Mz��7B[��,"��U��]�����ý� �+�O��Ȧ����\Tk��?�Q4>���SI�B���W�-�{�M�)t����Q�Wc~	8������=�+�\I$%�pbA�H���]�&�w�[L�Hx���D����
�,�й�q�Q qDA@�_���ѣ%�� 	\`]��$@A�7�
��|sLzK�Y5-!O������%���D<b���c�8�d��ײ��'Y��w��R"�12�az͋�n�E�8E���N�?V�Vgǥn|��<�sAM�Q�k�+�P�H(��������n�	l/fr�b͞�C���D��
��%���+.���S�l����Z�A[�B.�����)zK��>G��d��L<q_�8�n06j�~V?͘�r��R�a�Kc����5��{$�:m]��k*Q��7?�x���e�]ݰ��ձ�d���;�A\�wρE"�[F?���C�"��A{�ի�Y~�g�4�3�_�ԣ~���͡ֻ<�F�A;����D�у�3��3*��;Y�1�<��D�V���l���0 ��q�د�[�X�ļ�n�q����79�d�O�h]8n�	�<���lUuI�n�nE�I�$�/�X�N�>�ؗE.�w�sE�,!En��~^YDl�xm��cb���O�RTWt��w��(m6nml���|r||=E�A]_˟�ci�j{���xo!��w4�x�:�|�I��Ol��΋D����"��j���ȋ?����-�ad�rX�8��uuz��:iW�Tk�����_b����,����*8����ﷅ�˳�~)tW쥚u��|���-��B�iw���YR�H/�H�cF���v��M�0���{|�_)���/#M�ʰ2�S5Y��
�i�Xiz�Iĭ�Ѡ�#��K��?��y��7�9T��NRQ�����m���RO)D�
�:Ղo�klBK�<R�������F����d�q��~z���h���2*���,y���U ޑ�����)�@=y"����"YM���;_�-S�����8���*�)�z�+�HDB2�G=K�5G�w:��ԯgX`�,Kc��|���eK�rqZ�^n��B�7l}o�V`����CҠL��G�J� E����dj�eޘm�o�u���u���i���>�a�N`C+hr�����ȸ���6����o�Ĉu�$|���X�v��Ħ���\^�Dn�z�T�)�];mwhcU�X:�a�*�Qr��i�8��>A�`p(X��*:
�qZ}Y�yqcK���� ����Dx�"�1��o$�k�@H����y^=�*�o<��C�� H��cًrY�k��E&b$^�m��ۇ5e��@/�O��r��ɖ��
�����j
�������	݋�J�ψO'����������J}s�l�R!͹ض��L~7��;QG�&xO�C?�0I�K.Hb	�̴H��V�$s֨�����d�?�o%V{�d�6�34��oxek� :s�p�,�Gh�O�Z=��i�Pl:K�����AQu�Vjl�� k׹���:�A ���/�W��1��}��`�K����b��V.��$����6�C���<�ڂ�P��{WU��~�Ay��1X�o���Ԩ����TK4҂v�恿+�4���U_���"�p2b��`���3��I�P�5�KKC���KsN	⠴\�t^'��<���J������΢EcL�#Hl[�!qcq�K���2�K�K��F'o��Rw�T	��QEn����yQ�dhm���J���{�k�Z�qѱE��5�H�=f{<�4�7Xϋ����L���v%Fυ�DU.^�%�Ԏk�ZA��H9$!҂)�f>~�E��c�Y��K{���Q��|d��K�D�U�A� i�����ҐI'?(�} �v4�/*Mj�g���.���M�+�Qyh'w�\U�J��C���,{ﺔ�ӥ��"I�[�WX�翩<U���[u���Ӌ�����:��,ϳ�*�l�I �Y�+Emw����j�f�FP5��Խ�Ƨ�!wyR�l��E��&�.7b��k��Y_)��^�>0����������YP3��V)0bV���/j�K�I�ZiS��g[��}y����2~T�,V�JƁ��wZ�*�Xy��}@���t��(��i����� q��j�c�IE�Ų ��%ع��������˼��PI�+t R� �	rlE���C}EVWGJ�j���U~�OOϼ�XN�p�٣���4��(�]��f�?����{��8���̏W�j��� �-[��x�f�Uӹc�V]@`�%wZ����Rі�vj%V���۳�>N7��ݵ%&����쎒���]��5R����zP}b������;ex�f=�D�Ŏ�������i\vT�J�V
rG��v_����w�H��{J���l��a�k��䜏2n��Ë���zaX;ꮔ�!_?��b`��Rb٧Bl/Z��j;�n�����hjZ��J�Q�h�$���:�#D"o��j�>���j���ρ����6��{��/��q�l����V�l�)��
=:��-��g5)!=�pYvRyy�>I�+Q���E�N̋�?炦{�6sO\yg{=O*p�)S�VVJd�g�d�E�Q�|hu���^`�Jq�PF�SQ�e�q��=Hn��ǽ����&���Z��=��޵�7�)�<��Kp]�;�iR�8�L��<`�>�˥U�H�Ұ�a�k0	Rn�&U99EJ�n�gZ�!��F������(��>�ڱ��7z����1�3�<��]@��9����K��R+k���\L-����>����oCD�> ��ᇟl6�����WR-p~#vm�����������,�0�BFC���������%��'�N;}��_M�(v#�]�ۛ��T��"�1E6Y�W@v#JQ��_�C[R�qb�Uꤘ�'\��}��M@^����z���M�/��8w��k|ӥ�a�M���%��%7���H��͟��zu�� Yװ���#޿���ɝ=���+R �Q�zl�=�M&F���W�|;�V�����[	�~��޵�k�ͩ&��.�M���3o��e�k�vjվ��.�7�#��Pذ~\أ5S��իO��tS���5�C��]>\����{ �LH2P��d'&��)�F���מQTk���'�����w�ayF�uQ|��H��X��"�ޯk5�m;�u���|�~(Rdq���6�%�t�P��W.ۘ"��o�e�g�r9o�~�T��woޢ�ㄞ�$W��)^ _Er�,@Y>&��f�S�C�*�6�ql�k.�"=�0��\��n��0��A�u�'�K\:�c�uoPv���*շ��jk��x��i����6u��r��z�X�������]����4����H��y��mI��N�;ȟ��dr��[%0��/���Ɔvut2�q���p_�Rԅa � �g���w7�ˊ����<�-Kh�Ӭe�Nm�8��x����gF�,�Y�O�{-]�dbK�ԲF�����4�`6*G�1L�p�6�T�p���w��c����`��W�*�T�N�B H$L���C��)[G��\�����t����H���H:�v��K��6�o/y�M�b�R'�
����*Œo���!;2�{�ͤ���՟aY+�{蝌��m�|���+֧ʞf=���i!*�E��ljhvhc�u��[�P@��z��ΧV�U��;6}����u�O�UN�����e�(sE�54���\nI�f��#/~�f����^Ƽ�w��$�s������3N��`1+hꪠ����܈�+N�"��#���K.���TbAG�[�}Z.��bZ���RV{M��[��� ���-F���#�o�Q�!"����|l�؀� }i�\x|�A�*j�ƒU�ʎO�T�]V)�m2ަ���J�Eyٙ��K�FW�/k�l��R�ZQ�k�)u��c�[I���$e��J��^I�����_E��H��d�Ƥ����Ga+ MI���c�U��i���.�ϧ���V��)n$IO�dt݊cm\���Z��EE��&�M��	���C<�ip��4Ȕ @1�7���π�h�!<�$��-Υ�m�J�ߏcK/�J8��iTx�s�*6eW�kєQ#�ǀ��{SFK����4��L�A�}��9�b|j�'I����%Gl���n���}�s���ob�R�> 40~��&kh4��pr�r�+[k؄��~��k���'V�@��Ma����77��d��z�$IF��Dn���}�nV���L�Eh�[o�8E�n�  $=q�eR�;�wi1:��A5��3yO	!9���װ�p�����-|0�bS��k�K��m!�o%s�=��5��|�����;u�A�����\c����l��%."�A+(�d#�o볍p�g^�����^��8�&eV����73�79�Do��7��z���փ�܏��9�?����w��G�N�ש=�#�g���U��F|
�22���nu�p��G���R9R9Y�%O�H	��˼��C�fA�I��?o���T�߬4��juI��M�m1|���
�B�$ZHyX#*S�Wz��Y�ǌ�k�D�#�>SL*r|-��VZ�ek���n�8Cr�gMu-�q���bA���Z��)����j���v�����	�֊�+����u=�ǹ;��+8�@ޫ.%�����e;��{[�����1�g�~>�W��_P�M垶�o�j\vs�7J���c᳆p�q�^~_)�e���5�����Ì�^����w[>��1��V+?ل>w<�N�k���^���?:H	\{��'�cQm�@�7K鿬E��m����5��{�ߓ��ټ����46�[��'\��W}O�$`B6�wd��K������Lܵ:���jrհ�ص�3'������$����$��:,�b�G��J��XZ�6���]#�HU�Z�GO�PV��9�\{�A�å��qE�4)�2cf�����Pr��N�롯����9��
?3��c#B$(��H)w���'*�å�:���ӫ&��:����DZc�n�䭛&ց���L���WM?���f����YT���W��\���c��T�ܫ�@ �7�.�hr6��3�����#�ʯS1���{��]yd&3l>���EKm�ٴz9�E'����!`1������	���͸yy���z�i��qW4�}�Lw���� y���eUP�p#fT~�D۽5��mk�RE���wK9�V���w�}�B�N��?J�
��Z��JO�9���ޚr�i�)Ӯ��Eo�<�]8g���h�����S,��������S������F㕕�e�i�37�BK=��|��$��~�)�Sig|Ѥƫ����5��cy��8��������Ԓ�f��o�*����9/ֱ���;2���)��ٚ=�G5��}/��˄�ቿ�e${v�{F�z�Ȩ��$���\�qv=�Lj���F}��Z=�����k,q01V���xF䔨w�[�r��{SH�`.Z�"�]�7H�k4����b6}�,�{ʒZ�jL���]�]rU��iW��.�a\���TA�@r�ށ��:ta��A�'�Ľ��4�;���g�!Np�F;f�&R�^��Vi�̫�ϧ_��Mg�*�6U�FyC%Rn��bVK}z�?�}�{����E����El�$y ��z?�&,��}-5���^~�-O�DA��ŷ�jM��>��?��S_��q�X����ٷY#�L֝B������w{v�����z���m��pO��&�NEoKN��KT�B}�A���iw��i��|$(�!�m�4Z��6�h�;>���.\6i��6�`r��~.w��;�~#�V;_ŀ��\�q����;��)�T�<���*q�>-�ery'��������&5����WGE�}�
_E@D@I	ADZBB��R�v`�!U���FRJ��i@z��a��������޵��Ə�X�9g�s��g�g������I��/���o3>���i5�-� �M-��o1�H�Ӥ�i�387�#���h���y���1Zَε�`RfDgv�3�|n�Q�=���Uw̵X[W�+�UJ�ffg.��@a��U��*.��z'��
l��yb��GV�B�#�E�<��jbe%�\��c��L��u9�.�y�*`E?{�H��q�I�u���H7.c�1�O�A�/=�6��\��h��\ #�g�(A���5ў=�,�����E�O�U ���O�Ec�$��y���7V��i��6h���c�$/PH�΂r�J��!r�Q���r2L�u^?����B�����I	�k`�f��\�n�M�x-��P�\T�Ļ�L�G=tY[L�����68�6<������6}	/�/�<���W�V�?+��̵#9���a���'|��~DT�I��!>H��PƲ�@�ܳ!��ڒ�6�P��Q3��!�����dٹ���������%��Q�OF[;XLw?^/��p����YE���@]�(ϚZX�PQ]��Ǌ4��cD�J@E�"��W�8Ja�U��lz��i�Rq{�*��0p�B��-��X�6=^!�U��M��K��E-�o�j��qzI�?�8�vݝ!�������dB��X�)* 6�_S[�uݯ5�C�)�.�X/{��uf,b(�li`�����"Է�j��97\��+zh8��_��ܖ�V`s�u��x֯�m��WyD��kR�1�G����]b="Z��g�\؈~�6Ak:�a<�gR]�!�2��V@�;�Ř\��wӳ�S��ųq�� ���I��toX�3�e5��$5��mNUQ:_f�uM�c�6w�1�Mq$��3�U�Y�@v�~��?�����qj�����Y�	�ː!x���v�D�v���v�f/��B�>+��ϐZ9����Oٴkc}PF�&΢;.�oF��2k�q( ��[mL��=����|��*�<a���0��v�D��W�{�Ԩ@��;�n�9ܰ�AÏ��	ߧ��,�Ms�ݿOW���8I���{ ��t���ъ0�9S��F�d��q`(FS�*̙�<�H�'Z'��'��y��^�� ?�?[Ef�?��0]~1�-��Qqx��V�+��sˋ�e��2��͡&j�I�O��v�pcteq���9��(<���0v,b:��������4��^��iR�����/'![���i��(�|��O'q��3.����,ߋB^��n�䑠�u��ՙ�S߄�`�N3�O�1+B1's���c&���VLtW@�g@/�j��+ue HO�r��-J�*C��ÚU��Ȓ2��������-66�3�_kD^tQT,8مT0����֗�<k����5�/e���;�l=(#l����
_F�����������v�`W�W�;5��<�l�r7$��<f2�J�"��������Q��������ykM�A���])�M`�������Tt'Rz+��S�ZW��\=joX�������=܅R�~�I�N��:+k��Rf��Xy����k�L��Q����-W�\}
�C��-Z|0��os3ׁ��5���}��`��]V�iݪ�J�65���X W)��#9�В��d� P��a�����S0��=��<!:&����H8�y�Ə2j&Ԅסj��5��ç(��3��ypx9�����E�;|�0�ٵe�#���G;�ͳ����(�oZ����BkZ�����z1�m�NLN�x�r�֦�0��3��6/ߑQrGF� o�JmTL�ND��$s[`�X�*ێ��M_��K\��������F�f?�Gw�hK��y%�t!g�����,��l$�;:_!�d�h�ڝ���^\��4i��� 1�:��@�H��R��@���('�����[I����ϗ�D�m������ˋ�O��mq��\7����]s�@��rg>�.H9>���f4�@��&���!/S]�0֗���+�m����FgvW�kir����9s���C���f�I��I�id�>������T���8���L�ȼnf�Ԁ;b6,�K?6U��ae�}�y >����@&?N���(=X�TQS�`	�Z,Nu�� ���B7��Ɗ_m�t������GD��b5�vދ��v`��jnI�MB^�-�_A��I�%s���( @�p�C��:�����*-��8�] T�]�a�q��CK��ts��q���f.�*�#**|�-�P_8�4cኔ.^k�Kg��YkN�u���z	ږ��Y��K����/�g*?�N7Ǽ�CVI[���EPR{.�>I��oV���As-U��i�z��M��r��\���CkF��O/Xt��W�������b5>�
�S�,��W<�I'l���5�[7���>���)���ik��0�o��P7ۈ-�3���>�!b♷���u�Q��̰FUi��B-7�NX�*�eè�'JƧ�@���t]M.ҷ�4q�a19|/9��sD���hW��|�Q�޺����RŒ���G�A��G��̏�O좊��B�D�����&��bzP�8�A��şʾ���7��%����~����w�������@����&�t��b�=���vZ7�>�?<�X,w���<}��zt��J��?.��������!i��������#�(z��
���Ӫ#S�y�/h����}f�/���"�^j��mj��l"�f��D-x�G�^tU�gXǸ����"�_�:����ĳ71U�0����{�0g��^������r����徫�X�0��_���R�T�MW���5�yVsN(��9}yaǂ]C/<'`����m��˕��3�a�d�Y�]��)����O��@�a���Z��{�缡8��[�O�0">�L�N�D��T3��A�֚�Tn��5�I��"�\%�T6�Y@��+�Y�C-�"��������.Uo?�n���s��3���j�?�b(�-�q��&�5���ޘ��FXͶm��C�r��{����ꜼW�Q���O
�2�PB������|����s�3b�K�o���i&G�16Yk�e��,>ȑ�6*{�꤁0�ٽ��e����^@�B�>��ڇ䣀iv�P�g��"e�#?ؐ'���5�w<���gZ�hZ����`ҎޘHlE�������L����s4���"e���z�W��W�gѓr�Q�g�(�̧�=�HET8�زf#�Kpj���`��ј�������>�C�������a����-v(w�S���֝�	�����ΥN2�ϟF����,e���Q����M�y�(Ïm�8%.�G�O�}��(50������*�ӑ��쮹�]�tLًG��_�o`��r�%r�S?��v0��׮6(^�ۯk�E�7g�J6i�X\@�RֺP����,Ͱ,,Rk���r�����a/�Q,Ն�;G�tP9(5P��5�� ��xo��JY��;�;-Y|���N�3�X..T4�M��\�V$WD�X:���O���>�%�\�{{��
&�P}��;G'�wn]�1YG�U��U{p̗f|f�a��ہ�>�w@{f\p���p��{g����,�����cJ��`��)��$M�[���)s�kQ�sdI[nǏ�©FK޻�;!��EPNb�����x�{���/��D7��7�X��9	��Y����0|�4���`��y�S������ۮ6G�ܯ�Q������"�dA]�=l{�@]���e"����+d�@U�������v-�L�h۟��+��mZ:��;|V��b��y�?���';vTŏ�/�0XS�/3�;���.�ߦQ��d�V���4O��Z��i�MW�H9�U4hR;�ʫֱ�Y����U�	�}�]�Z��:4�0J���.���̇��43#׶��������� C�"�T ��e�̻�zғL77��uX�a�J�Z��W/��R5.#�?*7j��p�i�j_�b��Z�7g�g��=I��<"b����{s
x,^W�z��}绱,�;Wo���v|�iY��>}�@��	����4��dw���3�qV@���*��A�ٰ4��X�W��<��{aQ�n����Ͼ�nc�Ge��V�O��V�U��Mx��s�{s뫨O=�ɌȢ��E�ƾ�+֛�>����D�@=Y�5��F�]x��OJWU��W>�9��*�l�	��W�mIyLH��+Z ��/�թ���xVl�g���1�ͻ�CԩiCt5{����l,�-�$GS�,b��  ��n1�Gw��Y*����1Uj9���S�{rh{�{G�-���"�������	f:�!���!���������;����������m�<��i�F�SSC��B�a���0���1���cĜy�ӽ/�}���JX���B��ӣlh����Ej!O��G]�j��㖝�v��$���FK���h���,j`�y��JP���ww����"����BR#�ڵ�\��u.���q`���ˤF�
S�B���2q����wT���6��*\��C�.Zc"�}�_i����H6�&%î8uR^��eOl�?F(���G��ܢ�Mg!ﯞ/@�3h�K�й��R$� �Ǳݽ.�]xu���2/�᪱���e� qs�
�$M����E|!��)o�b`���=m�G�F_=��<ri���O�X�K���9ހd���c���1F.�!��u����@���6�1db�ߺb^�����U��k�O�C��Xjp�u��;�3_n�X>�k�3��s��<��+�5OӐS��g�^�-��N��(t�D��Ff/$b���X���0�8��*�/@{��)�79������3���Z�,Ǿ�kҵ��P?��5��JbG��xk>:�\�����.�v<w2%����Q(����Y|����5�B�A�F�{�����-+Xvh��лn��h(s�ZL5 |�]z����a�Y>�.�>�s���3}������U�x�@:������)��H�=A��V��U����h�F�5&�կ��{=�<L�����_ݎ��!�`h���~�7v
Ǽ�L�iS�"�~g�,���sC[���Àz��>�2�k3k��7%r����O]��i��� ��4R��.��n�]|X�bk�JY<{����R�^ЙO��E��"ɻ��V���Y��emB�,�ltkKDȬ~t�+���f�)�n
f�W�M�	8���q��V#	����F�7)���ӝJ��&	�א�:��E7	iOm&�A���8(����4_�[��J��Մ&�����N��� �1��+e2{~0���8'[ϴ2��4˲$˹yz㯍R�"`��+���ɘC��a|��"Y,���-���@@����===c���\݉LςI2��b�Omg�g7ݝG��3��8�;�`e�)���,y�_u7imZ�L+?��ۄ ����by�&�{��rM��Z���S��(CB��2L�AZ������oK�"@{K�:�ҾQ�:@;���8���{^��BZ ���-����oJ�ߺ"�	ӊm��
��k�iC�����3�k�B�`]�ˊ������Xޝ���U��9��?m����c�h$w�*�7MYF�5ϰ�΀�2Wn:H� �T�������2Gz?�ߣ~�j�Č����G�y��@��%���Tӝ?@%�4�� �Cr�c���#��	����nl=K��uwou��6�fB���=��*t��gy������I�	��N}�L�k��'M`!�,*7p�����^�N��O��K=f��c��)��M껆������6�^��=2>�㞺���+U�u*ew�z�$j|Եrܿ)G�qF���mf��ҍ�]�q[��8��	��u�t`��8Vyulx� �?�x��M�Ϩ>�N���9��5�O�Uؒ}��#6��)m?����ya��][�a1�u���Ӷ��cx�_�M�b]����^7���?�H7���9q�����{��o�#+���i���Qu҅���F�\�7��� ���z�1y�s~�js�4�*G�������������1�����"ϗ-��
|&�B��i���;�J蟩����~ '  �� ����������p�@~�1�d�ȩlr���@��b2wϠ���vGe�$�a��Û[�#�.��(���BiYI�x�Z�ި�nz���#� 
��IIK˭�*��n�kլ�LO���s'���(�	�ER�?_��9SUp���<�09VɍyY�\�NQ3E���;s�=<�J��6�,5������upt�Z1K�#��HϠ��z�l��j1����:�,�o �2�?:������df>�i5�;M�M��"Oګ5��͌��`�a ��*I�qP$$JTȲ�Z�[�B�B�7�xcw'�OalL�! �s��`,���z�@�:��G��C
PC��Kgt�X�A2�j�|���k�=��Ӭs�A�pU�P�
~���<��:t"3�y ?<P�[�U�W<��C�����M�u����bV�K�T,�b\+��!렝�N8�����6u��p�� ���&���De�&��_Y`�$#%)}� 
p���V��9�����8T��M�rY���g�v���W��Q�r��(�����1�Z�
�.�$bZ{�������O�٘J�=I)C��ǁ=A�� r�p����"��#}��p)�2�|=D5��i���|%��.I��j�<i؝���x��P0H����\�>�e��X�I��WI*�F�H�=�OL��*
L3'l�2����(���.��h|#-_t������/�{��u�"�5�]���`������=���������ߓs�~R�Lp:�^����8ȝ��f
��&6$�������P(}�(<�a:ԋ���<�-�^�z0X����C��)(d���^<�������_x1y	���z�tOy��w�_ݏ@�Hu<��)�������y���		<�n�����{ mۺ�^���;ϛ$��٘zu�)����d�zndD��m�+1!�؁�W	.�Hzi����S�i��R,���^��P1�pzZJR	����\��b]x�D���HL$@!�	�+����R�7!}�X�o�s���������H���j�~�[�m�j0�8:��L���㥟����{W�=�w�%���8;|��+��DE��Q���c_}�ΔQ�>��ߨ������^X��cx���MXV܇����f��Ⱥ|�b����Mh���X6���r�5}�/�!��a3,>a\��)=���e����3A6׽�6�ӣH�c��Wfɸ{��m0�\��������7�]a+-�l���*˻7����oll������
b^��^#��\e������X���cqy��J]�*s��[����0=�+�H�R�?F�7j�z�ZTr�(�>bh����3Z����4||a9����j/��b�&�xtO�H��=�'����!�[/1��z!?�,~�,xR��*ߊ�GF��X�'��4甍^m��J���tQ��x�t���L�pژK�=jw;N$��i�{se6�?�g�calޞ��l}�'ss��\�OEEƨ)�]�`�Hk���t�Z�6�$��9�uwSS�w3q� J�]�SǨ#�?e(F��r������z��'%�+|3�l^�2�k3����2ϡ�F�yG��Y�C�0_����*,] �b��aE����������~)G�-p�: ��A���[LP��1��ݯ�"7A�3U��б۞+�::Rx��Q�/��n}D1�j���,bݴ8���.��Zd��G�}c�&c9{�ρ���a�����԰�������vK�������6&�h\Xz�n #��*���\�I�t!-	BA���M����_/eu)N�"�����4�Q����}tv<�مX�0!�g�����<K�y=�I٣����jy0�q!
Jw���')(8��)�3q�PQ�N_V�C.h�yӛ���HK�����P�	}?����W���'�1T%��d��2
JJ�5gq���;��x�P�_re�VdnV�k�H�9�n��mO���gw�F!2q�^<.+K_,Nհ���c�>I��M<� �;6���������m�V��;`�Q��N+�d�0���5%����U�`�j���ۗHK����n��J�F@)�L��U=\��z��،���y�*����	P�t�ղ)�$%�`܂��;�$!��!`[KM�����kx8�R8�7JI*¸I�C�N�ZT�3���m&I��,���e��?4�7����@%�Tk/��N����!w�j�O��	"�-*"��/ �ډwV_�!b�}ɑ��#���gPG�j|e��|<sh�V_x4P�´���e�JR���m����!.���_���}$0�,e��kU��{U��ϊP3�^��\T���im��e(���M�!�\ʦ _t�Sd5'���N��T�� �E�K��jj�����S�|KT�n�E�'�D�rQ�y
�ڳb�7Y��Mu��
/�X�NI�(�`f���B]�	-[��D��zY'�Xm_`,	�̏v��;�����r�3���B�;�eS�q�:�D�~�\�([FX�>ԉQ�U����b(�G�G\���2�J��!�Bu80�U�*®IU��Qey���hA{���ʾ�ד��3��{�K<j��*ܭXm�%�U����1be�o�����z
hFă� Cޯ��3����JR�b��.vD��ϺPpk�J!����vn����1K��L7�bk�gY�	�P��Õ�2b���D�-��g�G�a���_��`��\��>b��x��b�5��H�B����Jz�zg2� XW��9�A�R�$�����x�v�8,�#g(�Ee-.I�_�D4^Y��
�9�� �����w���b�h�H��7R:�z_��jU��适Xo걪�E� ��pP�`�&5,ÖA��5�`k��9#YA�ɋG��*�9s�Z6񷇈�glo8��� ��؃Xm�;�6�z<?�Q-����g{_��2�
aԲ���ϲ��BRD�T�^��;�����K��Bf����K��Ǐ�0�R�kw�^�h�(S����1) ��{9�
�ڿZ��������ǭ��z�@�V��{��x���J��\�g��׊�t�d�.�<O���]�/O&j����z�t�0����Z6���n�ƿ�)� ���1$D˓�0�IA��C��^�N���7��i˪���R̵ͪ)דUW���s����(G�0��KO�����v;i�X��H�T��k�ZyD.�ynS���76ُ�j�~tٺS�@����p�;rb
~h&j�A���-̋�9���7�������w{�j���ƿ�j�_А�6y�$��\��d'��&|������1��4�«{�p�7���3�nJ6�^�l���\�v�忺^�W㿢q�qg~hh0:7^[c��i+�sM�(��7[������:p����"��(^v�c���⚿P��g>�`�{�?9��}������W�~��b�mapI��x���4��X��,Ql>��I�P��Pn�, �PӽƷ�����:Ѝ}�w|���L�5w�Hc8Ț8h^�Ie�x�.���SV�A�*�7冼��m� ��qy��n�KU���3���H��WTR!	9���ڵ�Q�F�ߡdP�S��<_����<��iS�[�8/{n��n�:5�\�R~"f��/z�~d��-�k�k��O�K:��L�r�k���5i�j���5eOeoN����h?e��S��1V���0�R�:�Ƕ[��y�|ڥm˺�I�yM��]i:�Բ��N�b#�����n�i@p�)qP�����TjP\�nU�F	I31���lU��)�hm��{����}�/VHώ��*�q����՘����x5��_7������'��;a�Q��1~XL���^u2� �8}�IS�M��;X�ժ�|!?�O�N[y�_ܘ)�A�������F&�9�i�1�ǂ��Xsێw�fs��^���E��k��ч�����
��ծJ,M��<��j���F��w��{���~2zo(���6}�=~�Ԟ�.b�y��,�,U�H�����9$�'�1Y�����%Ӱ�<�����0_	�$y���	?�(�_�MJ���㮒��%듟Z���3�"Ӓ���1@>e�%��_���.5ӎ�e��T�� �c�a��G=�
W�}��r�Q��Z�߹���+G����pq�B_W�e�2I�B���?U�jii��8�AA���:�P�Ǧ�iX:M�Bb�p<�G�>`�<s�0#���Q
��`�Z��MD+m$���"���'�?_�P��{FY>��ۤ]+�����t"�R�\S�z����7���A��� (Gb�uS݇�ľ/��T���v0`�ՙ�l��C�W�9c4�� ����{W&��+ɭ��Ȳ����yw$�i�~�W���N�a�����c�gE ��zX$~�36!X
uĽ3fN�3r׋z�����w��oi��T�\>��`b��)�77�70ԅ	~�1��Ζ�y��]�6��b��|���w�0M,��Z�������弼�O~7��q�p&��xkOq�d����c�T��:�b���_l���s7��I�c�V��VY��� @X��O0��?Ly�L�����]W�=���Ӷ�'V�A��#�o�8DEk����*��=+}An��_@�ϲ���~0����%����^5C��jGɠ?�6!����i��
C�.4.̸,wđ*Z�X';�J�O��f|�8�ryc��>���@��iRx�\m�Zz$��s���5l�0�wunk���{�3�����x�z��.�,A)��T�>���Q�I�)��?��b��㔐���0�m�~��t�F�Հ���@W^����(�w�x�qV�����D�\A)"�nF"#P	;��bρ=FM�;�=�^�?�p� ˧Q�G���dh�JQ���d2s6-z���q#9��}�r�i��ǽ�No/�=W�7TZ��ulԲ�%t�2:' $TEP���Řx'+�����d��sό/�ӱO��&<�@�I\�S��2f6�^��	����X��X�i��P�z��]i����4��&��E�PU|Ҷ�;Y��	w�=,�l�G�	��z�-�\��7H������g��!�[+�fU�I�z�i��w���T�ů����5{�2�7Y��jI�v2f8�1V�B���AJ�f����7�AM��ʀJ����{R�@������'@�l�,�L�=�p����B�Ѱ8��LV�x�k�$�U�W�g�b�[�$�өn��j��[�9�if��됬�﷘�ÖT��R��1��u|��1Vsa\S���.WvY���ͱ��k�nϿdk�Q�;_G��&VUa�۩4>w�Q�=��ߜ�S>W���m$Iz�	��3+�x�W�"���hD��fPc'O�� �)��[�Ap��DȡU�3��$�q�5J���Ck�_V�E���'m0d�nKi-͟<e��L�M�<����l1pL=��f�K���>�Lߚ߸|B�4��d��<F��.���=���ݻ��ˡv<��)��w&>o���_h4�bk[:��� ����O���T�:v�0��rJ!�'���J7�}ɰ#W��(�"�FY��eM�ִa`�}	p�������|�i�j���Z����X�xi�bA&Q��|��@�0�de5����C�4x�4t�o���\�-*�Q���@~�)��'<ܽ橝)���"��H�� 8��'G����ko� c�2�]��� K�7*�{�__�rW ]���XȣN��
�`�f��bW�;���m��	r���ܫ�VE��^-��>��j���n��3j��X����/�ݐV���2덫���)�y�ְ�Vr��2���|��V  ���D��EJ�U�M���ʈ�Ʌ�ڣtO>�7.~� 
ݐAo�}f��C�ܙ��&+ro������v���y���ck˩�sRW���c���s���&��$Aˤ,����W�ݏ��_c��/	^q9XX�ɯ=8�j&�l�D����]���/]�lע�#h`��XE�Ŀ<��c���t��pܝ���6U �'g�I9_`a��QVap�n��jJ�m�7{&�oo $���B�#O�E��d�Z6��;����J�[���6W(�b{ű����x�A�1>����� :�u2ǛLջ����y�N�S�wֈ8��ڃ@U�����Q���#��6g�r>E�u	ɿ��]��l�_�~����0F���/�zy������Zũ��{cB�	��K)�F�5��H��Xy#�h�\;xV�"�0��V\�O�A�z�J�":|��Ui�Iq�w	�г$�b� ��m�8'�G�?Y�?"�\��͈��yKj��,ZM���go��=%c�K��5�]��''���(ѥ�j$k�4������lːQϩ�673>@;R"��h��r��̠[?LU���ԋ�~e�q�^��˱����K�8��u���6�uj�f4�����г`�L�!�G�'�j�'����t�e�:��.!zb�*�F�|�r���?�}�A-�Y7��rK��QA����8�r�J~J�b昀��F���Zq�C�g�J �UhR�iMt�[7$��`-~�Aٔo��&�z��t����jjt�Q�iUA����&�)�t���S>C�����'��E��M+'s���"�!F�H��ۇs��<d��v.ҩ�+�(J&��LS5dG9_�;誠��J�-���v�W��Xo梨�;����x��Ix��w-���'{��	�m��p_{`,�Vlv��Z�/��J�&���+�� �7(���s��"�{���7	�{���x�{0EΏ#���E��y�l��4f����]��I�׃�қ�j�C��$�Ȝ�	����j��7� �J�ȡ����� ��Ƿ�9�"$�c5��9�X�y� �d	��d}B (o'ŚQ0��@u,$�ި
��~�Ҩ����^��Q}2j?yh �/����W�?^f�Q<��1��i`>�&� M3Nt �m�w1���
�	Ln�@0(l}n%�${�旤��*�X��W�:B̵L�h�l��r��6"m�︒ !���.뾺�}^6�'yB$��i���AoC����T3{;���j�4`�S�/���ʙִB��[JZ�L� �H�L��%�vѻ����~t o5"�^��!�!��n'�#�K�|췲bB����XjD������7az�+U�M=�?��] �L7�"���]}��,%ח �Ggs�P�������o?�ٟu(� ԛ_>NXO���S?��)����8b�N�뫤xG���o;i$�w��G<r�]����29L��<���P����z�9���Xi��C�ؚh�~�(ݱɢ��O`?5@�Y��n=d�Ϲ����:�x�|?��x��~��«�[^�9��F5(p6�^�dn"�����=�Ӛא�v�]�g��S��<�7'��ڝNW5D?,�ǋ�k9��Pn}aS.r�t�x7�vd�z��М�p��8�Aրl�C:p�c>���$~E�,u�l�i�3��Lf���~'�"��h�d5�Y��Ck`���A�I�ր��4���� '�����G�ݱ��C&��x �&�6I߫=�m�8�/0�l3ow�;��	�5S�5��5篽u��!�p�~ 8H��s��*F�V@�{�7Kq� Q�G����WIQ	��V��>5������n� ����������K���PR�Sf�.�'��E�T	���P�*:U��� �nAPr>RC���g_`r⭤����f]bL�E�B��t�\����<[C�N�F�����nI%(_Jf���-'Q��Hv+t���U��c9N�(�Ѭ<F��!��D�)�,z�$qQ�}��(l�H�����cr� �RS�V*Wx�� PK   ���X� ���� 
� /   images/38cb4f51-bc72-4d24-b782-e5d855ce8001.png�|gX[n�c��"D���  M����t)���!�H�.���*��@@�tB(�	�����{�ϛ�<<g�^�]k�k���*�2�etMQAV�R	���"�˅�_������>��B Ǘ�*@@ �o�/Q���&�#���sGM�׎�/�MA���|�6�&/ߚ��ڛŭIЁ@�@���\�W&\]L��{Tw��_����(���i�m���?t]l���c���c}y0�"r��n>�~�2�4�܇���y���:]=�*���u:�����,V�;S8ܘ��`��������Q�x�_���YL�F���N�I���[̪��9���?-�%O�I��;�rv(Y�J�ӣ��7ǉN9.]^;sn���g��/~���7��w�矤��2�Oߒ�~f�s���&�`O�V��2������[�
�β�G�~�z,�x�T\�Bgv=�@�(��5������ЅM�9���<�T)V��m���q�X�
k����8k~Y�֖���Q=�AٗmYo� "�~A!�����K���WS���>�7��eO�r�D�ơW!ԁ����F�{�v�ٺI��G��h0ՙ]8jY����o�/8�\����q*���⩛6�萕t��嶋�Q��E����Ma��?|)�?�晬BuGQ¡S�wf0�'����򇞨�����?�����}oy�{x*��h����,���B�4�*���caH���%u<�@�a��%���{��PZ|g�$Ӑv��+�>F
Z|�[\�U��5���:��Gac���|�{I�5�݁(������Y"��S�ʨ)^Q/��β��抖��h��/�Jq�U�_��:\�K��I��\�pk�*	(���t��Rj_k��i�z8-o6"���<7��f$Rv?��&hD�K�ean��AO������5[�U�tB��&�lb5�53$f��K_�S�j�nl�C[A ���>��fQ��b9���	Ysl��^�䟧E	���"]`i�ePybГ�O��ݛqo���XZ�GXP��؂�J_�]�Mq&(O���������O��oW��4����L���T$mW̄��-�-��w�
S���<��f��p��)k���N�j)����s��y&D Z��!��5�G�D#=�g��B�*�kb�^m{b�R����P�xs�s=����� ���R^�j��)���h+�ݰ����oF��3q���#��W�Ev?��b#�Ќ�C^�,�U�4����2��A<�z!�P"Aѓ]���~#)Pz�:q���Z�z����A��Un���@W4������AK�WI��=�5���r@�+J�:e/_��&iК@om��*�2h��w�0*��;7(�#"p��{�갥LƇ����	ý�b����W���ވ��DA�?)^�k�d�\X0��;0�FM2�%/�u���go���ܖ�Yo�� BH B$�2E��o;���v�_9z�To��yK�b�mFrv����f��J ̴(CN�w-�)�zܞ�1�i�Z�3�i����Jl�Y�@,�Q�=�kI9�N:[�9Y�CznE=��ܓk�k]��l�q]G<�����T�D�P��@�[�I�қ̺��e|�������k����dr��r@�B��S�VIr%Պ:���B`�(�i���W�t@x�Dp�o�) ��jN���j���#��A�qN�U�8�cE�n68�S���3b�A�
;yTr�}�Ȏp�W�H,�j�b�#g3��)��`F/��qYh��i�/sD�/��kF)�h�4gy]h8�����q�Y��Mh&�$/)�j�7K�zpb�;˥�6��Q;���S�1�G<�?���ϣ I�I�4��t7����bn��:�q����6nDrvn�8�LVW=�0i�i�~��|�n'W�x<*�L�-2	6�eDZ�k���
c�@2�sŧ���#	.�X��c�X�;J����t�df�� �OS�U+��'�f��N�atn�ɒ�o"���
��Ū�A���"q�O�7z���5�:V}�>̐0�RB�@�
g����ӊ`2�9����L�fk@�R�wђ��B�z�_�04n";،K�N~�g��M-����?�?��8�Zo��U�~o��*yȩ�ʪ�#!���$���|I0f�g��
��[��W��s��t��a�rє��p��ӂ���a���z��ꅖ=��'`%�������^��2�	Z�)XKS��DS��U���LF��A��S�å�X�W�3����H���_�\�+x6�xN�3n&؃Z����Nշ08O|g�����L֪J����/~[0Th�r��T[���1�1�)?򥨧�D�RA��S�o
_�!Lv,���zk�21 ���~J_"�&�f�=S���Sw'�^�}�����lbm�ec	��=/�גU��T&�BK���+�t7���l��W��͡���D���,c
&]�=-����xUV̒� ��K�ˑ&0Wn��Ǖ��s ���*��� �f�I�$/�+p�{�T%�U��O]�&�d���i�\�yꉭ�9�-��"Zg	�*��dU-���Eh��oe'v�N
_��}d��g]0��c.~�R���H4_?�1sD����\EA'䢬�d�X=9�� g|�|��FDt�Q���6�B.ҥ:�w����ZZETyVͬ8��;:�s	0��hЋ����x��Q����8IR��<�Vv{t��Y?$�f���<�/
7���V���!D ��S�~�J�g[^����e/77 ����~�9��-�p��%!D	ܥ� �	FaYAwo��-��J1D6�	v�C�Ӓ�~�GP�(�m����W��m�rsr�S7#�MF��������yyy�ɋ�FjM��FK9˭�M��w'-SL�7B��_�/�.�<#��eRHG�8�(;� *h�B|��5g?���(�3�ȇ�'�;�8�>k0K
�L��1zI0���،��D�S�,O=F�;����T��-�9Z��n�]St�#�AB2��'��)ν����(S%��T���3M��k�U݋�5b�~VT�����4��e<4*%�\�㟣&,t��ds�ψ�]-�V0�r�����o�� �����SIb��Z�w��d������e�oie��bA���G̴�7>�=m_1�Y�yN�x����C٫��߿B����&�gP�<x4�
��OIIi��4�Xwk��u �<�W�_����C�-s��L�����xݣ�J>ս;��Vxhhcס7��v�N��������Q��L�ɿ"��٠$3'gGp��V��F�&Nl�-i��2,x�|w?i�6��v&D��S�O!hm���$�/|N=ӗف�ޤ$3�88 !\R'�j̀�K �L�">Q+�ZZN����1c3t��\}�������oIf�ۚeeeFIǎ�^;C�����!Bx���|Uz��P!�������%�*�ԙl����_���b�Ť?������1K1��f�f"����]�8�{�$��YW�K�aM$����C:�i�%!Ġ����n����ү]hi�Bլ�uBe)����w�rg��A����k��nP���ve�4w�.0WCU:cZ8����S�������inW�7���u����R�ʢRPd"'�;������ѯn��,�~�`Lf*����Ò7���
�n�l\`�GG���x��7=T��'�W�睘�S�q�B�ʥ�4�_^�5�E7����Y���0}�;r�C/v?�cY�5ag\��a��R(-T�4�������I���[k~�ͮ�<����a��I��Qx�����W!Vf>�{�mk����VlX���f��iz�K��x�x�ʣ;*��x2�t�����OK�� �뮥���N~d6	S<P>>;�3��!i��gj�5`�L�8��p���/:$!y�Fx��U�
�V�T�ZUB��F�w]�^�9��D� �OAqf�`����kג�����XN���f�Su��wW������N�� �#���z�wR�s�f���KC�ڿ��M3���z*���e�I"B�	"B�f�,�Sb�,�jsxHa���rJ����ؼ�^Kq�8\��>0�0��
�:̦x��`|q-! $·!��̨DO���_�R	�{	9��eſq6��b��܀��w�q����Ԗ��{��r(���a� C���M�Bk��y��Q��T�Z[�l�0�*�l;M��ٕii~^(�HY��<����n�0 n��U���@M�6!��$�_{�#2�8Z󃺑2K����6�R-�S #�h��s׹��cNqJa�q��]�q��@�2�� 3�.�\!ݽW
����T��^l�����8::�2�]\����u*��L&>�;u�{��zX`�����P������Ͷ��x�;ف|�V$�@}�ڲMq,3ǥ�ӓ���<�t�f�TދU��{�Lu�6Z��Fl�щ�&y[��V�_]=?�+�
��v����p�i��{�+�M-�h�.j�{���}�9���bO���z`D*��
�6>p���҄���3����+k@M;Z̔+��E�4��J,6NP|J������H�_dѤM:���Í!�����w�QO�z�>[��OK���i-	鳜��m�!�!���Z0�L>�O���V�	neD����[��.��zM:��H��9���9��Ri1�a��"�Q�
�s��<.���"���CX'�觟��	e���#gjٞ�+)���S�b+�!������<�ċ�b��^���񇾢M�E& �]����5�4i-P���

�W;-�4�R����㴂�S��l=�+dvÚ���\s6��!����L% 4��[z&�����tL����3�9�x�n��Ά?*�ڣ{Ժ��m�d:���Sл<+|q�v�N���r�� �w99������5`@0��	���uf��[��޾'o�g-����J���tk�Gp�� -���w��㞊za�_ T B�YQU���1�������#b!�y�PT/�F�u�X�q)�O�:ء�٫���3��}���`�;Ƞ�=&�pyt�\�0T��:Sx�d5-�BTƫ����t$��C�W;H|�wX���qWXZ�9YwC#�%-��]�6�]j%�3_�a�tN�[�k����j��Uo������,��!`=I%і������j�%���72~P���!��s������䚏��6���gW?y�u��7�δ��·{��Sg�̺�׸�%���P��!6����:�$���I��e��#@��p�N-�Ly�$Bd���5e����bY�#�>m<G'CR�m#�g��c���������㽺}�G'�w�dkm���Kܤ�U$AK�n8���"w�[+�;y�3=k��(�W-0���� �#���oe{�$�z<38?��Lm���-	��NS����U��%?=;����D�Ϲ\,3�
�-@�Cf����
VŰ�`+�3-�g����Y�=Ʊt��2I&����1�)���v���[��
U�f�g����R��UK�vӝ�@B�߉���n�u���ȷF�O����$�e2u��i�E���|lu�̥��l��.B�q�
d��	�Hň�x��f�Q�6L/@��T�?�]�K d'�����M����7�Ĭ����g��Y�/��7҇�����N����Ú�S&��*6�!c�=�Sx���k��n3g>_AZK1��l�eee��R�Dg~��U`�Xw��P(Ɂ�˪ȍ����������ְZ�����
5�ڵƜ�Yjj�$	k���7��{\'����6�Lu�T����E�4�K&��r-{��B;�u9�{b���D�b�C�)!���sYw��Rpp�)Xጕh4u~�P��i��L����';Xv������.'vv��3j)��&�\�dL�����J�o�f�t���ʌe�p�f\+C�+R.^�(�B%�U9���KĨKgf�d0?�;�d%iD5g����x��vs>����|n�����L��ӕk���̀����!C��G>�
g�#O�o���y����H��ȺEp�{PA.�Q�`3�-��������[v5H�������9Q�Z.>��z~����J_�%A�!?�>ڨ��y|w������$6"�1C�r$c�|+��z0b-g�Mo_��ᴗ�o
��v��[�C���Y�[����u�'�HxWٿ*S{�e�){������L�Z+X� ��}��UF�s���J��[(�Q8"mӪ�x�x���D�K��*��������&d+o׮ɯ0�8�R�J�따��c!�4�8}?Ai�m�R�@���|y4'%��ج�'-�����7��ܙ��T���l���r�/�Sr��6K�h���-P�L����׏�x+�e�׺h�n����ߟ��_�ش��h���Ӫ�d66S��|�h���UWu;v�`�JEN6�zen?�>2�gP;��GI���j���X*1�\�w)�^���zJ�<m�;*�>�΃��!��j���St�L{x�LZ��i!�Al����x��	�r"��I9�D��^�V��O�r�)��5��e�c'���W�p,�WUcF�=� c@�	m9�`*�'��4����=���y��;�c8�[�;	p@ۇf�=���@�'���jԼ\�8�l����椯�F4�Xi��H[��2D���ɶ!m��W���2P�B�Ѷ�17v�����6orԵo®L,O�l|lTS��W���R^�~튁��bB�~�3U[$Q^���+Dw�!���P�)�nr�}�bJ��[y"wʵ_˫ ��&��uJ�i��h6񻑤�I2#=]���f����X�z[���h	i�s}�.������9��]΍���_���4^f�)���]��ݲ�azx�%����#��Tb�;x�ǜ�.�՞��<lc=�?9�9�$�Ͻ 5Gn;���ɭd�>aN+�Xf̼����x�"M�Vq3i�GRN�h�rg0��2Xs3N�-��A[H�M�e�Z�S��/Euh���H r��Q�ﱌ�ҺG���]���SXe>řU�;����9J���L ���Bg�+��c�9KwGtӍ�>��?�e2�2�"�@��L��]2F���3�|aO�r��$���T�N�C|�/Q�K�����E+�0�C[9�W�*1K/����匿A�B8�~v=���K��B=�r�����*l�"�K�3Y1�^A,��?�y�9��p������.ƅ�ac�-�|DmN}�8]�X:������q{�)x�v����v�ID��jh����!uO "ge�_�X!+�V)��a���㏺
��%��&��/��m���i�j�|�<�cFl^��cr4�vJ`��8�Kz�`�B1��׮54�[�� `��E���?�'������=��F)ͤhf8A*\u�jq�WR�˜;pȂI���Ս�BA�x<�N1�P!I�km��*M�6��D�8)e��U����K̂������~�vV�����:�4�\-���_��J�v�Y.�Spk���Yh��:~ퟠ��9���%x]�\o~W�	̊gW^��b���x���`T9���R~�q�W��)���Xx/���u7Gu�RP1��ؑ� �`�aG�������=Е5�Ѥ�	�'�=���v����d��߮Z�x��\�G��f�L�����֫ޯR�&�ʫ�M�`a�� �@��/���^��f��iv풽N�c�0G�U\�h�&����S%�G�`�M@���j�-oa�-�I$'7���ml�� 4��ɋD�w�`�׎�O������n�C
��~�,�WE�[;j~�d�۟\�r�ؚ�O(5�!���)��|dɇyti�V� �$f�p��
� Ɖ�WF�2V�L�����9֖tw����u�=���JK_� %��F�'�WF'�i�ǂ�/�$G"�N��ڝC9hAe���=A�/znQj{鷯T��$P}���Q��]���v�Gȫ��������0~�����.?�F&�v��
������ÞE�aM⋌}��@�җc��sW�h$h2Vn���g��ɇe�p@:_@�IV�]ܚ֩�<�TX���Zg�l��xU�7�-�����:��H�m��u�U��^	o�����^�D�dT��<Lt��_�8����͆�mKb/da~�@WA��[S7�N����J�x���#h����=��i?�~�@��m�]᫝��ߕ�<�,�����o��t_�k����$@��f�в2�0G��~���^�xnH�k�`���K��vO��rk&P��2��s��[�	+)u���c�"2Y�����.c�Õ��٩u���2�*(gj-��������O���cf��T��wN9i1���ŵ�Q���eH�^u��P�\>�z��!�><���R<$��M�vu�0R��Nt+Tp�v!���)��+2$m^;4J{�c�j3�C���j��Ĥ%p�)�;*��*n&����pOԮ6��lA�������=����ncG�E�٢G\�9[!!Æ��G/���N��<~,W��E�fșjqp��D1�u�������g���*˺ć�-��Mf����?	r���B��g�K�ea���1�Ty#�e�����_��o.�|�8��bg�(̅� �<���m�wvv�?:�ז����6��� �z2�51S���*7`�&�̼�BK���r�]��a�z��� Gm$*X�_S�zJ���6sҨ�f)F}��7/��-x��h^�+�:'����lA2��wb��ݞ�]|�M�9eß}&�u��w�G].�D��j|�4u/��y��_i�ߝ�;`ۃ�ڜ�II��zR�O�:��K^�UnT�:�������m�~�9\����$�ԕ��$"���p��Y(<[S뤓6���H�������w���yyIXwv�0X{��<2E���������jǉL	F7O%���*�Z�G��/�H��}�(���8�q�le��!�7ݣђ'�z�6 v�O�Hv�-\�����&���(�u= #�8�ࠗ�Čz�X��t{�$Q��E�[���`P_�^w}�h녕����s���҄CjF`�r���]�Mm�l�/,��9��B�iu�'�)v�7�\�+�����zqO|Su��u��B�`��L��ںك��Ml.;Nk��a�uϤe�=�~>��t5�Î�p�.�sqҥ>���<��h�����[ɂk=�R�:A9��FUņ�>$iE<��)�,_���IA^;�#��):���c��e`q�&�@j�.��'�&ar��Bi��[y�����s��+H���F��B�/�w����$t�K8g��L�����rW����۫��G���f�M�O^j����K�]o�S�_�o��ʭ����K�!�g<�E¶��Ⱦ�%�cr'��/ʯ*kE��G7���I�(#��2���l�|�Z�_VJ]�wt�V�W��T���;�LFH�<�U�(��i�z}۰�;��tir���fŽVQ}ݵ=��`QY,�g�M�W�̑Ά%�{��r@2@�r���&��6���)������؇����_Ժꍿ�b�n�b����9�H��W���W}�%��!�R7V��C���/@�������2y"�R��F�'��VŃ�t�3˟th�@����%���p�"#�b��o=��t��
K��fW��4ț��i��6Y6^#b�=p	;*:?�]�;C��]}�`mB���t�%ⳎS6l�F��%�Z*�5|�8��N�]��z�Y�o�\o������x�� ��b�U\�Z�w���3��K?���t����1d��E|�d4b�j�b�.���M2�1���8�<ha���^TU�/�
`�����#^�>ͣ8TX�*ג����K� �ێ,��/��$!Y�"I�!ʽB�Ъ���l%b�l%�Q����F)0%,����������- 13�7���|X1���^Ϯ����z���^I�=I�n�\��nU�2�~i����@@�VC�O~��&����@��0^d���w1�e�L=N-]��*?�0�ڪ7��艧c�"sT��'�a�wY�1a��^w����+��?(�G[��l%,�P��qmV���m�-��DWWך|���5�~/�՚���%9�Z���8҂��ۻĮ:K>�'Q�� ['(a�����������u��)�No���ɜ�
L�v]��ߔ���Z�K\?��@����q��U��۸�G�ѡ��.��;��rZc|��em��ж�1Q�R�O���u�؂�y�*W��Z��3�
aP�ڻbD�5����<:�_�G~;xϠ�e�ct�ϩ9�N��))��LA�mT�#��@�gW����xI�y�� ƂH9�U���}#�v6���שp��$���((�17ih8��B�E-����K_��,mVC	��
������k���.EA>�F�Kq1 wJ����\8�K3Bg��������p��|�'��j������ݣC�LGˤ��U����C�܀Yvd�����p�GO�L��y��,D%�UĊ3���쁼b����J�rL�--S��u<�t�=��m�{�v)^@�7��X�}0�z������hF"�Jkz϶��b*�N�]�X�������v���ݯ䇵j:]�b�0�L��h� �8���Id�����t��㒤6]��#���v,6������i�k�\�,}"h8��6a��d�k{�1��?t��������m���o������J��u�^YK����;���I��@2���I���>~��ΐ�*��^@�ˇ��
B Pd����Qypy*��Ip�j��6���7��t�r���Wx5�쑐}E���}@v���(XO���_�T�J[}_��Oz2h"HR@��.��>*ً� 7�Z��Z,	YK�$�2W`n���ɈJ�t�56���&I�B��]4�z����ᾭ�q�'vc��j����<7�T	+�=��^F(��s��i�p�pu��M ��w!�QC�%�{�(�ӏ5��Ǧ���%�-jĺ����~��>��J�;���=K�@^cč����I��g_�^���za	e�jwn��� �A�
�k�G�F]E�A�m��j�b��[e4��b��C�Οl���#���p(a�}g�$ ��6/���1�(mX�5��}����u�g��l�0�t��y��3Y�(o��|,`��������jqT�n�N��;�v�s�'�N#-���Q�m\͞�Im�]�ID��/�!P�{;��i�:�R3 ��������$Z-0�֯�X��Z���\�@��$z���u ;E�լ �m]M���F}bZ?LV�C=Ji�/�m�q���r�u���̈́���	*���0���
���4�?��j9�î�y�KU�2�uȗ��V,!�A��hxx[ʭ_ήqH�5�a
&q�ɇ���^������M'ܳ�}�T'�D�ԎI{&@������l/��G���a�WR�cPC���²N:�\�f�5��)e�n�\v[�ս�~�n_b}՛���W�Խ-��z-�}������`���3�"�J.m+4y惡����/`έ�@�D�
��X�B
��uԯ������)$ԅ��X�^w����#�<�I�Sꔾ��h� �B���)�.Qy"�F�Q���L�{t�ژ�G�]�I��`3stT�d�^�V�!�
�7��V��3��T�<<9
/��<LC�,��kr���'�Y��ܿ���ѕ��4B� ���,5΃@i��ūp-��bSh9�n���
�l�ԪNA�����2#9��e�M*����kX�n �2��`���nT䚽�c׸?��@&�QW�nǳ�Y��%]ʵV�=�4��ٕ\�k{�`M�o"o:x8�0y�eg�پ�2��Y��`�5/kMŒ&���B��p�?�sN!J"ꎐ��=Q���9O��]��s):�IB����\P܃67cU�E~gk��Ӛ+V�ϿdCK�+iTYl4���Aԅ�І�]:��}����+���㈆y		4��R���^�T����ǖ�d�Q-F����������3$�\��o�j-���.��\W�D%9�u�4x�n �ݰ��Rxtչ����E�� M�#L����R@d�B�r�k��5���J�2�OY�`M;#����#?!�o�x]�_��:2�@יv���ܓ�__E����v��[��E�O��2���z�܄��0\V��Mk�άap�9h�-_���c��m��F&�yl1K�XMIL���kuV� �rJ3���G�R8�YZ�m�< E�F��K}7�X|��af#�W�i��Z�Ɋ�/6� wsf���w�kP�W�Q�f��0�9��=���h�eH��Q~�%�����ǵ>�7�Ӽg-�<��BB�.G|:y{�޶���p\��P"�d��~Z�,�z��ե#E/V����s�v�M�5D��"o�N��a�;v��}����~3S�n���{�X
[�Æ}_eu����Vy���.����TH>�=��r.��t�ut��W~(bX	p���|S�u�FH/iL�/��a��-��?�E�eY��&���d֎��Y@��a�K�0��{�uF��Y�����R����2���H0]/�c���*6���	̴�������������n M�2�O3߄��Bl�2�n��k\��vp�-z�~_�>)*����)��I��[��'�߷軧x�?�y���g/���wMVA�v]2Èg*u��.����6F���3�W����+$j�mWrR�[	gpq	�F߹�O]�[м�"K~8�|�.�:c?M�]J�9-<��7�R�kZ���l����DK����s��1��佴�*��v�ϲ�8�1�ͅ�g� -���<����7�2f\�هQk�F�M֡F�U��F�S*
P�d��I�V��|�J��i返���@�ؐ+f��^#1&4%�;�ŝۛ��1@a1k�vV�G�b��݉�wGR�>F�F\h,���R,�>F 1����ja�����o����͜��0��D�&��0������6Y!j[�dP�#�sV[)��i���`�x�b�����P�Xr\�/��谖��G��3|5�_��{QONn�, �K�d�+�˶�M�)��L�7��b�S1?~��@�o	����m�ҷf] ���J�o����H|�19\x�ڜ��5_���*��IQSS[�~\���W��)��Q�������o���I��O�*��R\T����E٨\Z;	;��3q	��*��q��Xѩ��xB�x�>�sq�B��o��}��{N��+I<��#�+s ~wz;�>�����T1�~��bf������کj���ZC?���^���j�.������	��S0O���G��*��\]u]�U�MJ 36=���IK���Y��a�Sj�Ϙ@�L��	��Q��7�'���Θ�"���l�� D��(n����3RY�����l=S�%7�k���X���2L�@��X%�;"��"$l?��0d��
$V�۲��t���\�V���yTlo�%D����� ��D����m��R��!lg���lz�����}��U���>�	�9W��.����<��� P3�g������Z�a�*J�F���n�K���gq�m�aX�����T�����c���4W����j+_��I��#���x�6w彣�����W�c�m��ū��<ϰ㬨�t�\;��W����@�r*�
2������#Zؔ��[���Ԧ^B^��[�V����Wq����N}�I˛��d:)Ǭ������RD/-��6T;��p�ro�nsm$YE(@AD��ob���ͺ�`[��ؗ�& c/!0(4����f�&	,E 	)�{y�X���	3�OU}����`�V$vGtjk[�[�.�Q�s��B�MhL*��W�pr*���3�k���𯆀���;�\�y�����_f�Y�3l&@���_+d齎-H��3�2q�iA����q�]�9J�V��#�@�r�\��DjuݑV���WZ�[�b�$g��J�I���aO2��<��F�||�I#�T�Z;�x�����`�zP3Y/����1b��D��;��&�dC��9�W�<�V�󍾆ZH�w��ƨ��<I�~��,)��Ҍ�8%:[+5<�g�6�u��5_8��)::��Q� ����?D������C��m���]��s�^�^k2�@�-�i���$��x�g��CB�U@(��29�W��;�;o4q�V�m��$�y��i{�ٻ�����{s�YCm�'�5&�7�)�;6���L$6�ܑ�����d��UH��'�A�Z,���n��iF�ݖ'��|)��`�x�$*�u�?__��x�'�n��Wq`��$�(��Cxk�<�\�6�������w���O�Ņ�e�ЙyL&�>�3_��� t�.w�g(���z�-z ��>c)q�}��YL��ǏN�P����U���Ɏ�[5�5H�d����j���0F�Hw��xRb\��6`R����h�����m,���d�a���7�t�؎qCn���e��=�b˵ä 2�BU��[7�"p��g�'S��zo0}W���eI'�LS,�Zܻ����8������A��p�#�|.f�2���ñ�r��5�u9�3}�M���3�|���X��̵��n�Zv��g(ǔ�]͚K;��V{2.(��F���镵��%�0�nR���LǕ�a�H����=*�V�?9y�������?�a{r#*�:�!��'J���H�А����׌T@�y��
����ٛ�<�Y\'����-�F]�r�?i��~�?A0�/��멡�!���KW��t��d�K-�o�Ʊ���Ά��lSQ�k��n�E�I�J�BB���:|�^��=� �D��J%H�S�(�Y�*p�Hfq��`��z��{��n�Yl�MT</<|��I����5dt��ﰇu/^*B��Dnǚ��[T���p�,n�koP�
��[�Q8D�����p-�qV��vyO�}����v��E���o�
��S@a�;���[�3Ln]�p1�Y�Yt|��[�7
�����ɤXI`�w�Ĝ�#_���tb1 ����|�NU�Rp���9�qo�����O����E�D�+��!�?�ޒ|<Ϡ*�d�dm�#��!���-y�\�?ފ�F4�S���&e.������D|G�Ą�M ���S����Ы�����{d	��a
O�����	��F�Yy���@aA���k�9�m\F�KW���z�%#)����9�R�XF�^l��t�E�����Tm��d�|���@7qЭ���U2�A��u����2O.�mNտϔ9�v��U�q"֊(��Ξ��/�[� �"��ٴc�"�Ȼ��t��� 1�l�bs���/\9��kN��BH�%���.�J2�\��i�q!�4/*y���W`��]j����_��>{��pd����g�+���tC_�Em��X�W��&uAA�W���ɓwR,��R����L�R!�)cQV�| ���$�] ��T4xo粰j?�����݅3ʕ�Yǩz?����.�ru��$�=����]r�ѸGmPl�b�*�f
fN/�v*�#��m��Sx�\�p���3uL��$jkA%���ע�� ���;+�wA�V� �<�=hU!oX�EF�;�2|8���	J&�������yL�a4����wE8�N9�B�2G�@8�<�Ը���u���/�z7 � �4�Y�&��{i�b�B�|�XN�cÑ�	��^�	�g��F�tJ^�
�ѹٱ�Z����[�Q6��>2.�od�����,W�r�{�C�����t��:5OO.����_R�ޝ��x�޳<��D�S~�9��AJ㺷w#^	|�P�ՠ���<)�E�H���x�S^�2�v�b��lW/�V��rK������E�u's�d�_��eٵ\����4-����x��Q�	�һ�C�C�{�"����S�Ao�����<O�3�]o�-��w���7�r;.$2�O`W�A�-H���������-?���"�#��	W���8楙�̉{����OyQ�Rn\�����4o���5�j�b3zu����u�D�9���PEa�b�2�3C��Jjb�^7�|w�/�(S��de�$�{�^c=Pg�Q��c�ys��I� G`��\y�9����3�\g�%�^T��ܫ ��u!}� 0��37�=0���p2m�~+��n-1��KT��=�a'�FP\-�v�pZi1��pt����j����7�b���������"����x���j_��!h(]��3O�D�F�O��f������{7;(8�w���ȍ�����'� ����Fr�&�H�����#��k�=2��rb3�����|���G������]:f��0Z�)�-ve�2��*Y�ŐCѾt���b��f.�/rk��}lN�]�Ȱ�l�˻�2I�wi��z&c :x�H2eW^x�+���p���.���.�_K��������ۋ0��|��}��
��u���>�)1����/�QO��@w*�Aު����Fd~7BV�4�گ����*=�6�Ƹ"^x��ǻ2w{���{���r/���m�W�9��ӎ�[�G�Ӭ�Po5 �����Q^;,�<�;�7#j�$�#�Ck���L��r��[F� ��Q��.��z������j# ����� ��DRnw�k'N�F �'�UA��.>���.Øn��eo^�ɓi`Fm��?�o�Hw��&� ��~��y���:8�V|N
�d�ȯӲao����}�&e�Q���]!�5@�[@Ω��"��b%���}K��Y>��˿�`�[�2�9�2Yh�I�W�"�Dޓ_%�5(y�<�޿�"���k���H���j�0��e�V�[q�&�ʣ���k��T�JL����q���X���gUd6�uGj@�W�{�0穡-�������t�Ɲ���ُb�p�֤tDѼ�},�J��nT�6��Y˂�<=D����ً�4�"`��a>�ǔ�T䢀v��ϼ���6���FQC�o ��_�L�<����F,���O����) �y��y[ R���C�=��[���W8=�VE����W�5�vac *e!�� ����n&��c�0T�{���ݠ"  9z��c�t���=����}�|�����\��+@��}�	�،�� ������9�V��������/,��i
/-9�̚�������sMhL��QR?i�2"���<�e��>���;�/�VH��,E�U�c^�ΫA�.��W��O��ԩg�F[�{[�xVh�`Y�>
�]�����%��GXk�]�2�//�~{�S
	�{]$x�e�X�|��y���^��!����oa��˹�	�^�?e��5ݰ5x��|���ʹ#WS�\jU�p�i�"�=�"⺎v�`Q�N|0/u�ad�}j���/�l�~�HBm�bu��n��&� ����lo�� r�+�	��w�_\��IS�e�z>�A�֖ B_$P[ڠ ��@�6J��|uc����?�5X?���X!�$��˚I�l��AM���k�)3y_�#l��{[v׸;Ao3f��;;��ٶ��|�^IPs1�\͓�H��k\�Z�cU���[��!��4��lqB�_�� ��P������;��Ϸ�j���ګ6_���[�_�(g���A[�vKVl��Nz��g(�릋Lm���%����bD�I����g=YsL#�\�,�l=ȱ����J������6�9��ܣ,������sq�r &`� ��4+��\ӳ�F�q2��U��m\���B�۟?��r~�dKW�jBb�Qj��򃶻��tr�I�WT@@JL�|>ب?\#�{�X��6? n�F�$��f;��� ��������d�����=�{�#OWv4��D	"���γ��nG� à�6��o��3���=F�$3��\��[/��	_�U:��Ơ`���G��9K۔'a���#=�=xA���j�eJ��~� :���&��+�=�����'�W"��Y����Qx��Vٗ�<�o@�rO���@��$`����c��L������v,f�o�>���":�}y@��m�����癁m!4nD�je�4�O<�����PN����e��B5�z?!�d,TSdwHNV���pF�Q�{���t���u9��a;΃:���X��RR]S�\��A �?{u��2��{�������\e���wx)���:��5��HH�xC}U<W⻗#˶; ��[|,�����9ZȔH�r���������X;0����R���7��;��9�e$d��>��ޡ����o�c9���& XP?G��9�H��bqt���3=/�2�[N�3.G��Cl�w4O��8���"G�5^�]<[�#���9����֤`�a�/�����t���彔��°u���ް��(,����鬵���1�7�3�j��,��~δ�:��R˕r�(��J���\�ǈ��v3��/K��a����FN�w�χ��:�{-L������!f�srC�֪�ߕZ	Tگ��7�O���~�Ё
n�Л����� ����?KI���1S0l.Lt=@��Y�� �QF�?]��E㺦��n����t�v�nxn'�-�y������"�|���w^;�GGof�g�f��3�Ys�ٹvv���l���dL�d@��5�aIپb�_m�wg�`:i[�}� h���Yv�5����zx���Y ��l�Pf䦦���ݥ�Rx����{���s��sn�}��rc��yO���}�hs�S�E���%W�ўOv	�H��,�4����{{9�X�{)/G�g9����amQ�иe�{�Æ����Ꮃ�v�ߏU�D9�J�^�Hdl��B�8��ˀ@$k������b��5]a������O(���q�T	�i�vLIiI��T	s�T_;�
��~�|e;K~�!$��d���s�������s��.��y.���zAe�M7�=T՛�O��~�����
w�f���ɨ{^3R2�+��
+�	��I	"JZP����9��rg���2����mN��3JՋ/�n�g���5��GT�0}�п\&�"��8׈	�;�E8�f�Oq;��^���
A\��]pq���^c��σ	��/�̖���Om��2u>�oT�_���v� ���)]�p���nn>M['�� !��!+�l^��ъy#�~Y~��gw(j��8
��I����!f?$���\aÏ�*�ru
�vvV*щ��Q���0PPK��CʭO��P���K�w�Ú�� ��-�Z��G>j���	�)+�������Cju:�	��aA"�l7�^Z*"���V��w',c���b���_�:�������U��n���˻��N�k'h|/�G�\�F�"�2��!9��O����*"\;�'��eh��ؚ�GE�X���W��r��;�VW�UlUZbt�dEbQ9n����{��R>�_�
�#ٱ��'�	��؆_��gpG�ǯG��'G��:j��cj���4R���I��'c�J �K�>��Mٝ���j��y�I�e�7o�b%�K+r��.�n�4���9̘~����иE<�[��ą?��Bs>;�A���(�#��ݧ��!O�����-@g�d�Bn����4��H�;-]�{�������=��� Λ��E�F�8�aOާŰ����v��#�ꗃ��]Zc�:�k4�P�a�Ms����VC�����S*'+g������x�b_�l��������pFP�]/	:d�-x�F>g��!E������1A(/��Ѡ���#�L��A6�թ���ڼρ��wD�S�� Wԍ)Vf�Pܢ*��[��v�R3���������6u�#�V:�o?��P@�j��!��j�՟�5�7	�ڴL���<�!J.r&���|\�y�	�'g�vhu�R,��K��g�kN������J��J�d�Y�.��/��;z�w`t�b���R��`�P�E
�]l��9�Ӂq탮�,����*!�'�� �O������!�C�Y��(�m���q�����	��"f�_��L
d�Ch�����g{�oVV��"�0��z!����i��;5������&r�զy�OTy�d��b'zuc8�:�<Rc�F�A�A�j�4~����9*��[��VH�N#L��j(�MӽM��K�rm�Ӏ�Ms=��|��DF�)&�"��ϕi�6
6�E`
f��[��R/�D�մ2DI��ߪ�db�������;6�ލw���.vdaS:d�P+|	��YɃF��R�cO�4��9&)��4)��v����7�	?7�JR���>PNy�O1�[�^nog�ɷ��t%� $}n;��{��(\B�҈n��8`Y=1�۟㝡Wa�MO5_����]��2Z�w�������`��\�Ʊ�鐑�a�i�J��0���$��N~t��g>"��~�����T1a�h��}\�4�S�>�������3r�m��*�OA&_�iq>x!g���%Q/�u�ؔ�Cx��a%�����ira�2.YAS^�U�l�?���V[�'�~|����F�C�����,մ�U�W�7s��>���{Mi��5Z�:�=}��m�0���莙��ߊ�Y�e�6D���әq���ݩ]A1�e��i�e����&=��lmn�5�KU�3.��8O�2�' cU'����oU?l�G9��!��Y�D/Rs�ot�N�y��۟���^�6��L&ߨ�֋���YG���ˀ+�{��9ޅ����O���,�|D!����˥�^�~�Qn�)*��\�CY�8O�/\ԃ)K2 �����1_�R����g���7�����\��M�vZ�JJ��j߷��
������x�@�W�٢G�����*��{h5#%�fͫ���&!���;�0��{��T���F�Jځ��qp�ßc�&M[�k�Ӎ�0Cvy*�I&&�u�_�m�'�ήW����������buJ�}�D�Vݶ+9�A�En@��y�:]T��DXE̻�RFj:!Xt�4����z��|aGC�������
w*��t�N����$���ɜ��f̶��� �O�j�-����rSE��oc|`�9[� �?���v�*�Ѳ݁�6���Z"x%����߳ T����"_���|��9L��a_i�e�Z�&e�aXUq�8[�p�����M�z�-Q�䔪g�go���j`�Q4����������oh��t���w�Fv0�����3���tHu�)�$]��"�\�m{�Ź^_='F��R}(�A��et�J^��)��oW꿘4)�@��q6G�[��ʮ�&�	���o*;m�V،%�^�iB�o��y)�1@l]v |'8��gs�����{�;5e���ea�!$��Tb�t�b?aF��W3�V�]D$���R2f��x�Ú�ml���������>�T"2.�����Hc�$D����}��
�z���l�k�@%�����a�,3���D/�x�|=D���&nڋi�:6Ǧt�Ҋ?[-j����ۖb�'�2���	�]塳;��}�;��:'�k�L��!�[�
��$��>�?�_�=�ٌ�;����ML,>�����1�|�W^�KN�	��+��e�
�E/�̀$�3$�*�y��׋��9ާI�g߸:���������r=2�a�oe'm�g$�t]C/Ul�h��48/��T�>����d���$�(�y�yvQk~ş=��2A���v c��?��?�j�O �:Z�ތ�:	�s4�Fl��q�����G�>*��Ns���7�v\څƵ++h��J;�'��wΆil�_I�O{e�MĊ�Kr�6�����#���^L��g�&���,e_��b�%o&F{9�z��O��+�a̰�q�}�r	�������~��/)\˒���ɞ�Ϛya�n����񭰍m��}��)\����%�&����a��g�w|��\�)�L���;w���z��|Ϻ����n@�ȺՏ�fvzҳX����V�CI��=Z̠��)Si�$�W	C�ɿ�?`�ۘ��.s({ob ���c����E�����m���w0��@�;�@k�x$ָ"�Xa�i�R,ee<0>��%�l|�yw
B�s�Z�=|���W�Pۉ��Y��ɿ�3L����3ū��N������vP���'����6�kT���uYeM��O�K_�ޕVn@>�z�uMc�)V�38_�N��t�Y�.F�p1��
#kbފ���{�-����x���>vw�H� $���QU�T4��>�����x^-���?&／nЭ�� ��&6j����S���\�������d�<�F~������4��e�����9��ƐC�奴�]�AJ�|��nۑ*��}�_�S�K�X0oYV%�35���&lJ8\�J�݁�w}Ao��
L�� ]����u�fx�o�P☺�����j��44�@ڕ4٧ݩ"�3૦8F˧>��E�|��� \��V����+�*5\mٸ�o�fg�`R�}}���B*0���+�O��n�pN��e��rb@��u����KgT�} �o􎊀Y�E�l���es���I��)]6�P�PY6�SxS���L��Л�����o~�x1��O<@�{��ߥ���"}1LJhB����"z�#�c� 
�{�|�e��uh��e\�FA��O,�n�=�?��ܵ阬!_�mtn$��.�QDuX��B�j+�o�{O�Ǚh�V���(�V��b�b��K�p&�J�5g�
��(.Gϝ�,�]e�� \�v"N��[g\כq��G���2�
��+�U�o�b�����ة�a��S���Gϓ�ZA�K}B�A�lw��Lp{k" ��@ᭆ�I��f��C�
H���ˠ��'ֆ����IܶwIF�@V�����6<c��7:�������(�������:����Gg�Oܓ/��ɶ��cb�h|��x�>r����Փb��+e�P����#�d�i��=?�s�(�v��]������o������h����W�z�t��P�`Q_�����/�޼�#�wl��*���5N��f*�RA���c��\Yo�3U�q��U�(hY����յ]z���1�
���&�+��ԃ�#"}�i���Wl۾u�s���[t�{�5�8W���)7����J����΄kjǩ�%R����Zi���j�%*��f��y��?)�n��:)=�]�>e䤫��.�N���1V�=�x�t�i�2�)�S4�04x�hԾ��`?�XoNG-�Tݍ)�����V���ՊnC�#�V��ķܼEk
�0��q����xF�U&�H���N��u [f��zK_G�Z�ڮy�zEd0#U�Z֠�K�oe	�f��lr�����9��@�;�k���1qL{��FL���������g���#.�Y��2������g# p )�&U�ht�t�ns� ���wِ�+�٧�o�j��!)�l���G�F�>��o[�+RQQɔ�hj���hw�Ym@t������޺g�}���qZ��
N��7b��O�Z�������,�FXW:J6�AB'�{���j�@p��}�U7_�.�U���Y��^�p~��5����`�#�nm^�J�\�\�^K�B�zs(�����w��K���yJ��>=��ʅ����
:��m���N��:o��Iz�"B�b\.{,٪7ҽ��w�\�	���5����tQ�Ȫ̬�+M��0\�'�TE��[��M�-��~R����9�2V��$�\w�nq���q�v>�����y˪zz��K_�]�g��'S�̶�M�NJ�3��4� �ͪ�OR�Tͬ�����L�Y�W�a�e�M��֔W������Z$���
�
����O�/b�]��\����77�JL|�\q(y�Q���K���t�V�6�Ě,L�{���T�M��M;���.�	qsJ�"��O�9���^�|D���oט��<c�|��t܍�I��8>�h�U�U����uLl7��ѓ��3i��E�C@�qC��7y%TнmO�f|�}��K���lƮ�	��DDQS�&� 
����v�R�5�~���)�bu�������T���'?���9��~�#��į��/}f�@:�-did�[8�.!����]G����߱(����Ր�(�>�I������EO�h�lI+�fz�T��K�V�?}j�ZJ�� ��{E�b��ӈ]L�����ֱ݈3w��N�u���h���V�,	�H�b˼�-d�gHe%�l%�)ò׈���������E��L�cJW��U��K
s�tlygggtor�?��XNDAl����F'���_���|�A-c�c�;T�k�p��J057'0��מ^�����qF4�n����Z�gx��,�ƲQ�bSvH�r	/o2~-��t��%�>dӹ��i�����^�b1��*�v���VӔx�\���d Ӂ�������$�'lm}c��saIT9DL�	h�*�77�#q�����r��-GS�����N�z�n����3�����1�v�E�G�sU������(����w�5G���{o�����^{X�ܷ`�MOΩ���$ w�Nx��wI�egI�T白�+	�P���u��<ʋ�x�1���VV,b�r��wtX��0<��G������^_S�af)��Y�<�����E_`^��J��6@��v�k4��,�F^���n���� �?��mCEA�2�N45Vc]�%���N�Q�*&3K��?3��������>��1�(}���n*�6*�c!����t�\e��k���D��^2����=Y�t���"�oRVO�CB�p�����l�����*�V9���^Ot�̪Kq��7C[�OF�D)˳��*:�E���cRߘ�
+ɝ���>�hxN�Io�?�L�p��'�硂X��N ����T~o�s��&��ț���)M^kȰd�i��W������ޯ��W&�X�yi�sy)L�.a�Y�պ�;m|'p5��"*G��4�޴-"�K�q"�����a����W�X�SU)F���������(Ժ�u�@��6�/�$yZ��_J=|1M�qp��Ūz�����^-G]���8A���V(�� /Y���*��N�����ʲ�Z�_Q�1��"w������E-��ŲgW�A4a�ّ�se"���[cK!.��m��Uv�~�eֶӮ׈-ߣn<_�Ԋ�}�w�&�Z��ƘVޞǜ�l�n��l��.�H$���|Ԍ��6q_h����g��Ɲc:
+���\�aE�Sxfu�����w��i��Y����3dy��@ ��ly�n^��ai"#�6��}����N�d��!]2i:�ĭ*�ng��醇�:N�,igrfr,���u?oʹ�������=�85m��P����o,hZ^Ӵ@ӫ<��4����=�`���_�Ϧ������O��1Ѯ�꾘ir�����\��O����ߖu֨����i����_}�3تbFg�ɏ���/2ɨ�� �C7����xiz���o�3���[����Y�6����Uq��)�U /0;4��m�O/�..�L��b�6
>R
f�}1M����q�=FHsj��'Dt�͛A��`�3��������z���9���H�C���)�� (�6�B���m��ھ4R9~�M�ylO�h�6���4lh��ms)��Tm�z�I�$�}�G�0������A�Ұ�br�I�4�/�wvj�5Zxly��?�=n�E�Qj�8��~�g&%�8���SOI����,j�/��Դ�M�k��h���t6r	{��?T/�կ�/k(i�V|4�t���qx���4���a��X�/[�ko�
����C݊���!�����x8����A?�{�y��y�� ���^�G��d6T|�f��c�����pt��;���j�07'��C���٢i�Į�Wv��QC�٪	�c�W�͉i���I!�}e2�{+�EL���B<Z�j�e��]L�^�,��zw�:ܽk�cZ�%�핮-'������[�h�n�SuCnB�o�j>֑s����،�Rv[U�����>�V�b��-/,y�?Ø�z��f羥a^�rÙM;�/5��W�Ж�	<�>f-9a�~v.��&,�Es� W��1�������x< ��&�)F�P����i�*N"���p��<�\BB�n��p �ԮaM��w�cf��&���4���=>��?O�V�T)��A� ����;@�DN1�kF��Ʉ��$���� 6 /vH��G�V�;�����s�;g]Q����L��w]� kW	�Q�D4& ���`]�Ԗ��=��t;��έ�y_�~�ݺ��c���c_���hY0�K�"���H�Elʝu�c��z���#}b:+H�/C�?��a�r}W	��>U��݄�jS����|�"�~��|�?t�{��E�����q��u��t��|fUZ�Tσ��u~'����^ x��\�@2K�������+ ������n�8>�|�dP��:��f9ejX�

Sܭ�U(�j���͛�Q��G��M����&�#��.��]5���['��$,�_�a�I�F$�����۫�c�XWM���Y�j�1��"��K�.�^���@X�߽�C/27��kc9�l:��e�s��(��P3���{�}��٣���g?Q�
'U��1�m��\�{6�ҕ7�=P��:�N�51ǪX:O���Ku���%Y�츍\ ,�:r��5H�iJ`\_z;\ޫ�H(+����s&I
y�(����q��{��r���SS<�K��TS���?c]�ö�zWPLW��B�x�J���8�$vs�}=q\�1ӛ��g։��m�5�.r?d(���}���x�/^�ԕ,�.{��_���b`�q�����a�J��8A�����mk�`���7Uɋ�a �Ș��a��l9�=w~ϙI_�#�I6���뭬j�"5���z�5Z��ZWY�@�d �Ķ���7ih�%�"2H�#`����C@�9�=�nm��v�4�F'��̙[|��>vB�xM�f��&
�t�<1>�rHl���Ŝ�������m��FgKp�~�"Zm��{�l�-v�e�}��/%���n�H�s�I�~HuR=��ӷi>@g�^As�^*��	*ϟ���	b8��/�fVw<�e��=�b��z �����ķE@ߟ�**n�e�ZNLVҿX�ݷ� r{ ة���H%��씌0�^���E�����У�%׿�Wڰ�:-���l�����Y����h
�4r_N����ϛ[����ʋ#�;Х���<�F�.�ܜ�OM�]E��[���}y��TP����Ĳ�9�K�_	="R5ap���R��&���y�qi��Y��n/��F��у�s��G0��Dye�e�[��TMqd[���V���+��D<-@\��(��Id�&N��.�B��j��]ʚ����-cs=��Mn�i[?�o�Mȷ۱2a�\y������rJ�^���3���m��AQ["򗂧��?��A�T�T���{�S�0�Ŋժ�w�啠X�Wv�Q�wZ�r�Ne-�b0���!W�����?;}lmfc15��o����Lѯ6�"���`<��VT]��L}M��T*���4�w�_~������.��Cֽ���1�R�nndU�G�0�1'�i.x�Y�*��~._�hW=��.�=�P�ˢ�;���E��8ܑx�A6�V А�	��{x��4����>g4�	�]\.-�\{��Dɭ�
�=�D�;N(��ڞ���B=��+5�����ީ�_��*b���iG��Wl���D�z-2�d�>`H�$�#!)�!4vQQ����������oܘu0�p��B'�4���4+U��w?X��6�����|g~�|�����g	����w��kI�(��q��i%�b���D��q��O5�U�%��0%��Xqu���-زq�61����O5-�fi����k��'�P��g'�ce�׃.�S;eI3�MO�f�g�����n�i����p�SRmj%O-G4�������Zhc{�>j0���D��e�rѦ�v��9��Dp��
Mo��yO�WF��#6�j(Six[�����M��׼��$� �*{�UPI�l�@_lw��[�5\BD�8�A��h�֐@;un�~�.�C ��@(!.	�	E�.v��e.64W���.QQ�-��\�0�O�Ą��|��Y�gFS�4���d_>��	�E���v�D���N�q�?k��ɱ��K�]O&6������D���<
�L�٣��.[�������c~À}U$���e�C��#�z�j�)�M� �6��~	|���'l}2^%v�zRҮ��Y��?9�#z�7^�P#r�J��ޯ_��:���s��?
�X�'�j�Z;`9����+���Tl�m��Nf�����ax��K���>��1�n�)���L�A-/���,��l��, Jf�z��{�"���jTe���fKZ�~��q�2�_i���R��}�4�'����"PPX}�O*4��x���T���H���DnF���~'n�B���A���� F�e����C�	Ա�6���
�~>���rF�٧P'Hמh�qs��W1*����[�������w�0�}N؟�C�|{ҥ�ŏ�[Y�[���gz%U�꥘��z�$�T�f�:�ɗF%8�cVɔ���`y��ٱG�[�{CkUش��'���ɟ{�1'��mJ1��9aͪ��B�Ͱ�"M��zI��4�Ų�v5�+}>�`X��d��M���8W^49b�Ӫ���p��Z����U��ۣ�5�Ϋ~��g{$����'s�S��
�r�ʵ����1��})�K�K���Ʈ �Q�ROX$��ʿgC6��ٶ��i�3�l��O��7���=X0jQ_Ѡ�����MUx6�����|���X&^H́7�
�L��D�Mr���V[�QX��
b7�5.df�kU����M�S?�X�'�G�t旲J���gR�3�>WO1�Q�szȘ��u��-�J?�ke�)��?ԗé�?3:��IIQYNwH�H����������������U#�5�K���]h>���#<i�Y�"�S�d�5�,����7:��AF��ӓ�^�����p�m���fYj���Kϣ�+�C5>��jW��պb%��/EOic�.�R�B[A5���3���
3b����ձgKB��r!G�����<u���.�]I���W���jE�k�._X�`�3�H���IL�B��b.��*�B��A�O1ș��~�vc��p�̏�-l�$�Ke�e_�jR�#Y��\l槬H�4�צ|�#��[#5��Q������4�&��(f-�\d;WੌY�Q�Q<n��Mml�+)���p��u�|h�[٫A�x�@��DٿX2''��ӓ�f2���_N-��`㕟��*��[,���=9h��C��J���F��:P0�M�����������`�@B�S��@}ųFܗ@�JX��o����%T�%
�8nI����.�J�9O���&��cփ[�;g��\�7�au�����&kb��U�����`���D�&�P|�NL��Р��C,���e]�*���.�5[������v
���}���lmR�͛vR�X�"V���u�;�IB��/%<���.�_O�(
w=�LyU���Ù�\<W[�1�	���&���#�&E���ĉ���N�s2��-�1Q�`�Y� ����pi�V�G
�z����r�mte;��вԍ@���V��SUwᏦn+��s�{q$w~�o
���u��A2��֧��Y�^Н��)�"W�6M���W3�X�u�i`����Ŕ�%�����\qlX��P���YhFV[:�s4��.� o�nv'��iy'�8��Np����ɧ�<�����<� ���w#$Ď���D�y��+�+�["�8<�>b*ğ��UΜϟ��(���2
��i���bwr
�m`���c�}�2��
2����@銕:m��C,�g3�{{u�����q,1t������I��"�h7��̺���_Q*��6��c*g�oȵ��i�(�V���۵�A�gx<K|����ܶq����N�������\�ӭ��W~P���2b�A�Щ���b��ѷ�&��(�Ri���5j'뻝�����JT�z#�, ����;
��p4Փ�r�|5�7� ")�C��K�H�PNt�l슦�z�
hB�����o
Ym ��V��]�^�x��_��l��&�x&E�l�j�$����{��k��G���z��������%�\&�T����;j���������?6����fRN�Q��S1G�1oq"�ĲX;	a��_(2�Vd�<ۍ�Ze�?A�}�\7�}��lH�iG����QD��X�yFG�K�ǀB ��BЗ�����S���h�WK�_t �C��!���G�E��ޖJ�O��o{�������z^�Kc�4"KfI����������H!��b�m��ub@�jh�&��Y�ڕ���-�����{�޸�]{$�H�@��`<�
��T��͌|ۘ�}�i������]�q�R��p������F��\C�����LB�ȚܔZ"�B�#�ƃ^�Iܨ*/��SE���r$g��f�M��F�mMD0y9��$�݁�OJw�� �#���*��.������
�՚5d�;w�I�7| ���`qj�$�܌q[�%��Bt�?��*,�"a<��^����5g������<�ug%r]
����Ҧ���z�l�nl���Z�Ը35���Xl�����[.i왙�f3�� ��˾9u���>(3���1�ٍT(Tء�T�s���oSB�~�ӊ����Ѥ]��΍�=,//���3+�F3��9o6-���w�{�����]/��K2�����܇L�7�A	�x��I�K%ץ�1\]�D�H�&-��*����O0+nl�"4����1f"2ۦ׳3˵������M����[ٯ[���_�+����]}�B�y��!x�c :����
6���-9��aY<GR!*2��q���e�E��Vc�Q^9�?B��w�4��mȥ���!�tu�<�U�[��Wײ�_]Ӆn#x���0:Kã�r��i���[��+��癔�0�=HUs�E�	QP�ӹ��E(���^d��D�iU����k�{�� {�?i�|ÊP���a��yZa��4)�#m2˱��ƉMk.���־�Z�<N�{LꞱ/��,/����X]�[�,��/�6`���'C�|al�_��=������D���@;��C��i�!´s���t@�����mJJ.�׼�bz%^�YNg�t�����9#H��G��(�)��(y�S�ӿ;o�yQ�[ Kba�*�8���5�����\����O�3,�kP�-F���1v����ܕ��4��K�=����$���iNK����+%v���n4���+۔䜄������f�{~��J�!I>��d�=�M��'�^�e�yx�Nu����<���1�_C�����}��956**�����~{g���v�m�¨��Ն`��ZO���ىD"������
~Mq�n�q޳�o�`
��S܂�'�->�y�%�L��_5�3�����>##C�)��R�Ѳ�>:&f4��Cِ�"�&�z���b�pggg>Hc0��ʋ/X?���6�����_i���������0��0�p%�w �v���C.����?<�������W����ꥩi���x.~��]���3���\�-����F�U��X0��^W����r]P���G.<S��ݙ(нqd�PO�K���"�"��+gv�����w1		0���D
�f��.IvEf�$��#��{�������J��ûFϟ�W^dLv�q5�QRZ*�
��Y����7��,0bk�0Le��FGg��)�0�lwr��v���.�wFrE�E�M� ��0�G��;���y[��1���+�c��+�44\��p�h�3[A��aj_�z�V���Bz��57��~�6�c�	�>55o߿�Hy��B�"���K�[\6�i/�������`'��U��E� �?�Q��ty�4W����{,R��'�ˢxg ����{���	�JJ��������V�����bӀ;�_C%����rT��#ݾY(e�؎A^ߍH�B�|
��[4���A�R^\5H����!�s�=�̔�����w3��W�.%��OY<���6LNA��u�,!�[p-���?ن�U�t�D�w|g���Or�[���ڲU�^�N+h8���hg�/��<a�ׯ�������E��[m�.�?	��A�� ��ۈ��y��?9麿!g�EWR�f�c�	X<)Ĭ-��t�h���V����rz����0�/Lth	Wwo��A1>��s�䉡�&&�������-)��0N%=�|o}�Ts��{[�H7�)����o"R꯲>���Z���Cn���y���z-�DEG�B��^}#���H�,A��Yv�;�ۤ�
ȕ�A��̕�HM��
��ͤ��O�A�
\�n7��H
����$u��K���$a0o��c���c��U/�8�c ����[��H"�ߘ.{��N�Ĝ��J�e��ћX|b�}g2��:�_�tZ����7�}r�2�C�~v7o��Y�����	��s���Ň�zol�,�Z�q}RȆ�5��W�/ffd:7t����l	���kx�Myw�N�&�w�����I�_A�\����a�V�S�߯)���%Z~kM�5��p6�6CF��ޕ���.��//+��ɑ�m���)�˫Y[#����k� ����c{w7�|HF#����BX>���A2���5'Ǉщ�}eu�
��y8� ���, �?k)(|������r����505�p��Z�b��}8$!�k��1yR ���z�� � ��^5g��V��/�eZ����' ����]]��	I�l��81lׯX5����@s�����,ׯ@|����'?܂.� ���C";���7��b�D��������A���e��6X�<������~'��g[k��ش8�r<������Vz�-O�dhg�����r�30�0Ը�?3H������}�z,��pRDꐈ
�!{S�<^��'N!�ۃ�8� #/�F��F �X桦��Pڋ/�ZZ�iоT���:��`�����ɏTփyz
rr��1����5q#�- �d9���v� �^=C�er$w�_%�ڈ҇ư�1)�,�D��n�~�l�p۬Z���E�"�+e?�̷J F̊����Qں(X�S,���g3kyy��^�_f�ANEe�h�V�^�v��h���}���5L!1��d��I]A�W��^r�* "����G���}�x �]7;�]����b���ؾ�X΁~�� ��g���Y��ׯ�h�J�D�������9���	o�a1�?�����A�o� [��E� �w�c�Q��{?���sm��/�YV������XE -Z��8�@r���l��V�ENN���Q#�|��*���ÂժirsssB�P��,V��Q+�{��\�	���l�qq)��[��9ޟ�/Ԙ��L`i_���;ޏ)dcg�R >�0�z�6� A��P�O~<ow(����U�D�0bJ�ޖ�`jH�����ףȘ�lŞ�+���2~�zlp5���	�Z�0eK�z/0f֝r���|������@�^��߼�]�_�K�H<F��nJ���纒s�P����%(� ;*���5��{����3��i�ͽ�=\����ht��v�F��|�{�,��z�������%������#KK��W%	$D��i����ז��,�s�:�mJ�����c��C��z׏(�<�����#D��Bo�<8����;Z����&�R���֎p.�W>d�KF��t >��zf�*#0��G�T$� l�~y{{d��v�oi ��5Rj���G ������c���aQ.�������(�$�$-��H���>hdYn����sT��l��dm��j'\'i 6�ع�U���ө��7i�L��3/�0����j4Nn�w����.@��0�ȩ����
�a#����˭�Z�r��O�����rG�u���iw)Rk�3,!���a <�)i]q�-�+�������r,͸ދ�g<�Iq+s$C��i4�ߟ�h_#��g��t���!��l���@�R�i�P��K@�Y:�U���Υsa)i���XB��77��}}�_~v��{��\�9gf�����ة����힄��㽒c���<}Za���+u=k^H@ ,����L�ww�u��h�=PkdL
�[5j�����0iTE"1e���CzI��� ��������)�4����;��x��h���fhm]1�Dշ%���i�1�z9kk�4������?%Zɱ��Q�6��g������x�#J��Q]�z���r'E�WLO0?)�w��Y%��2K�,HB��\�4Da0[7[ί$�DGG#7��f�w������_�Խ��b��࿷�3���	0Μ���oP'	;�U��ăΊs��Q;fq
���+����^���n��Ӝ٫歟��d�D�:[˂�X��o�����Y�P����	֮{�zc��U��� z���"�]ޞz|`N'�%��������Kos�z��kKat����q�����#��3�N���1��#ݜ��7�>{�1aL�7n�|>豴 ?��bhC�\YuJ��&9|�����m�zC	:Q��h,�ڧH@D�m'>�)5�#	\�04,�}o�-��������[�33���1s㞫b4�� FDW��}F*-kg��p(��ID����<��-3��V����{�m�Zl�#f���f�}C�v�P]G���K ���\�ǖ���3�+..U)/&	/ہ�$��4D�������\�:�#/e�m��ҷr`d�ʔ%r�F�B#hK�����Y�}�8���;�ش�2��p�Q���������A]� �p�.װ�vGeJ2���i+x�U��SZ��F�jt�Z*ae�׋��`n|o,��S��(%Y�����A$�ra�y(c�Ĕ"����}vM�����#�mm.��(C����	��Ŕ�Ə�$U�uYRJF
�5Z���=�A��w@<��
�`�<)��<ĘGg�C����V����}:[��6PSS�V�T�S���7��"��3�����mqyy�ؤ��ֲva�d�n�՞��!���e;z��ׂ�.:�+�s�I�2���eѴ�
W;�E�o���L�_~��*r,ߙ�	��]I¼�0�f��~�$R�SY�-Z���&�"x<\i�֛��0Mf��&��P�����n�9Z�
�1�@��QQdk�U^^�>�� �d�Z��8�?l���
2���]r��nn��եN
��O��G���a�_��'b��Π{s���8�P9�ta��i�DQ�E���/��y��uy$b�X��8p]eX��|`����\*&�3�ܖ�Q^M�vg,7Y�p��QA�Q�^Ȑ�_ߐ[Q	�{�0L�?$Bُ���ގ1u�ӹ�e:�7b��Ɨ������)흩}��nP�.�'���rd�b+�o'�r�"0��ZaU H��WX���D�����9p��^�^��T[�����HĔ?1�s�j�f�JW��򋺭���%��qI�h%Q���#��M��$��?�^6�j�,Q}U�9��t+Q�����$P1�ۜ;�;�Ő]}?s��O�UV����x�_���bg�m�w�#�s�����J��$���w�.\�r�֦qΛNu����(湥=&n��z����ꨞ�^�����d����Bb�O�^5�����}����{�.a�TV�cي+�����\7�'pڍ_\��N90���?�w�_翍��w&?��*��z=W�~�L�f�{YKS3a�q��'�GG�O��gp߀�/㜆��g���������9���x+�.�4)G�K&�z��b�A���$����x�4���D����7~KK֦ff�)d�$+��۶��{*


��4yUw�ڙ�$ZH�AZk�q�������.�7�#��`i�=:���q�c�]�K��W�T���ފ������,9g�w�g���y�q;��K��cȝ1�kso�؀���U��3e�c:g�f:c1Q�7�w�BF�&����������<�Tq�n���¥<����l6����jQ�B ���hhdo�����>;� l��T�Xd��m���k�hLv�d�s���W[�F�6]�����{Ƕ6sU�@�C�?��F�N�h����kL���&�O`q���{t��k>����U�5I�\��2��-p(C���Z�gנ�����ڜ``��g#��x�@3��UlհU}��Z+��ԂYt�(%��Q-+0Ԙ\Ԛ��V��㫊N���ߌ���xwN�^P�K2�����g4����C�$��5}�PhtAFƃ��׮���[���.�7���z���9���a򡆺�<��(�-o!���gYQi�SA�e\tI��q���� ��!���g�ZG���V��sS(�Ew�Ы�{��2����y���򋋻s��_�1�geee�@����J||�����Q���P���*��Ά��7J B
�C�G*0t�r�tS������ƽ<g�䟓�jM�7u���5z�����X�܊M�t�R�P����"�I����;�%(8Xع�Dw���B���X��+�184��O��*���%b\��A4�L�0�%�t63'a.����8�K%��ƿ���lsF1��(� �R���[�3ZzX�c��Lr����+η��~�9G�e&�Q%k����,a%O������տ�`���\�����}}��������,&�����Y�;��%��߾6�L�5k��5Z^X�W���@��<X��H|Τ[�{� ���J�LXWt鬝��#�Hn��{���/��8h�$	<��<7����͎��3� g(��41�趴��~j��M�2a���E���\�PA��ٮ��$�n�/��&<1}ڴ�#'Ɣ���3�tb�1�7o��<o�f������e
SM���̏~����H�������� Ԕ���1%S(,4�^ef�ۊk��A�/�x�
��q����3�����\�CSZ3��/t�z4��Z?����8��c��sk�NJ��kOGG��YYپ��Έx{A������rOr�'<�9��r�j��ovM�c����F p�!54����.p�&�?;r��?_+��$�䶓SS�=Օo�Y2��4;+��v�``�g�}�ll� ��(`������=qrZ���XQQP����R�yYY#YU���b�g^\Z�hY 3O�ɇ;�yg!�Q|�a1����m6�.9�_'��C
��걸a nL���m~�}�R�/V? $$�oH��@��#�1��������(+K>�P322�-9�|}��D���]�u�\h�^jjju���}��i�Z>�o�P�CdsP�
��|Z***$�.�3��S4�/�̸�I^~���:����ꊒ�}��g/ ��V"��ɞ����t;�KX��3��_=��^��Y�]���pxT�y
�Z�ݫ0���	C!5�������gd�;�q����M��R�r�7�&��ݫd�#Co�"����7�Q�ۍ�ʗDƯ����CWV��Y?O#��u�fkO��W����n��d>R ������Z��,�Ç�̓�
�6Nt,�ā}�:�sF=����e�,�6٪�cj�ι�=�{*f�ך�7�?AP <��V�\���9����X�%s%#�}����W�wy�Dp4觊G]�իtn��&������b���1��-��"V5�&pv��l�P���6�r�� ���9KH�;,��`�=������r��oO��yq��CMU�����6���в���%��2_9J���K����F��~�A a�2��>�I�G��G��s��B��m�V#����bn9�ua�~��&?���$��۱21	E���lk�$d�U�_:
ḣv��x���b���喳�(х.�Uh+�D�hz�o<�b�g � ���yc����[�b�2�O>��a�^__���a<�]�x��a>����|��?��&}����i���R�_7hY�1&��?�@���8^�[]A�x�����X�Evv���Oo�iv�P�Xr_{���K�+���K��Z�a�s�N1�P��;�M�3���v]�r=�}���*����3��u���߀���.]��nh�*	����}x`��]U��{�@�CUE g�e�2.K�� �~��9���4�����X��������,���c�_�����ME�"�#�A�讟S�[q?�{��㖗�V��n7T��2>�**�r,�!vvv^؍755�F311��׏�t����OӸ㔇�@�cp��s�
����*�`�0מ��>����Ci�c����H�d�RF����ş���݋�>�fn�Z�u�Gu��R/:WY���::��:�O��n������^ K�1�D����	R���R�M>޽۶žG�Լf!�er�P	;fEDD���/?��s���XvCJ�J˝�0<���jt,��o�G#2?r�jR�R�!p�_�v�@�4q���{�l�����K�]e����Zʚ�J,�0����>����0�^��1�<�	M?�>>ޛ���(q�m憬����q���w(F�ٹ�m���s],,-��J �� �!bz�D�c!۶�=��p��T�#�Hל�;�L�K�,?�L,&���A��ϟv������
ŝh+]�S+x7�U��2s's�������k�m/�C�iY*����֟�c�{1�$!Y����Yl���0��5��d�og����� �zř����W�"�P�l�ߏ���T.$��7ꗠ4Uh[;�N;����+%�tg��s^�5K/�_���DϞ�;�E��_���`H�h���Uuu�j��x��["�98������L�۠����O�C'�<�x&~�}����S ��g]�:�4CЫ�ߚ�m���+��\�u{]�������Ko(D�'�������1�!�5���TZN=�}��K�/ķ6�r�J�0��7�i�D��ت�=�������e_��7(��$�ZR�W��u���&(<�t|�z��`m�QV��_/�a�d�9#��tɋ�6��Ŷ�"�����iR<Iʌ��A��5�\�bҁ/��� ,��w��m��6����|�`=C	߾)@�K����I�\��J�^�7J��+�\�z�����Fd��S��~��/ᆊ*�~||E
�����3#qq�ٹ��qm)���O����:nW ��ӗ�A�|���{�Sx���Z�t]�
e�<�0�G�{R(��ϜI(��[���jTB�A�!O%3*&f֕Ik	[��l��/(Y�������G1yihj��s�4>���F�����5�ϥ6������Ľ�(������H̥��\ۀ�y�	��^���PJ��:7-��.æ��۰�N�
�P��XCZ�m9.��#�X0��Qm�u�d���D��PS3.��<����A���z�>���W.�JNl��J�Ґ�n��1V�&���^����������LG'���]Z�+@|-�5���FG����.q��L�u����uYwfn�s�e��#���&`~�{�ɢ�I_DDu���m$����EE.��ő�`�U������.k�G�����gDm���R���|§˶t���c~����N�ފ_�\2Ov���u�IPǘ��cs1�a�m��7���ޠ���x�Ժ�H?Ҝ�\=�ma��}�3:.΢ �3N�^\���0)�ۯ��V��Ýw�E�1�n��xxE�������GP�n��:>����)m�6�QM3�2o�b��Ś��o������af!9�����e� p�F���5$.�a�N3����c���<��ɓC��{�%���#�1�p�b��T�a��XD[��,�x��5�Jԏ�t)Z�'�'��ј�������F�PTl,�+�_qHCCc�=+[>4 �Ɏ_�b�Z��������l���|��U/ў����Ӂ61~͙��K*k}? ������|7�1�*RsOP�����m|���5��_�,�ju��8������b�a��Bn���mѨ/��=�6 ��?|�xF��^�.A�j��ՙ�vr^���X4��~u��V��7Ԝ+*�A)\�E�|��'�l�E�u�Z��*�ÿ��|^�,XD��촶�����ڱ�I�Rg��Z}Iy��}Z���\5�+Ub��D��z$ե'��ӡ�P�$��S,z�wV���By�e^�Q�N�U �lF*U���܎w���������p�=ru�˃9�4���ޛ�����8�O(���m��KM^�eJ��{�l9�m��ûq��$�z�$���zRl
��XX���n�+M�>j�v�5չ�׮\�D�5H��� �
-H�e�|��ł5d�B��6�ￂr$������ؖF�%Q����Y�0��d'�՛��N��y�{�k>sQR��1����UwO>E[i=|�N���P��I@�\o}X����7�t���J̕��C2��Z�5C��*'�O�eee"G;S�蹹9A\����!~Y:�Ҩ��ş��r�Q�~'Joi`dgr�υw汹��M������ ��?���	 �kB�6Xiܷu��a���3OOo�1�uŀKoc��w?;ڜ�i��������M>\�~��0�B�P	.��`�Ք�[,��4�@�i�(�kdh�(u�}�q���ӽ7��i��G\��C� �T}�U�][�h��4���QQ��ͭ�e�]%��k�C2�v�S�4׭!+x&�S\�@�s��ԯ�A5e�>�������Ju Q6C¢�K�»C �@Ã��x��&�&F��^�OtE�}��x�����=��?�M[厦MOf��וּ ���ck<�ا`��PYZZB��Z9e{��cwfh=G�`�����k/��,}t�?π��� ��]'���i2��.�j+���e��<�l�r1���n�Б6n�Ⱦdx�t�xҵ�BO��?�����o��\\�Um��E�/)�^�V�
XR�'GGF{./WTٍ���-y{�n1ݝg/���h֧��cvv�Nq���kp�^�cv��X�'�� �y�`�}?�V�b;k���Z':���Z�'b7�٧b�e���a�Ϊ��Μc#�����+*B�ٔt~��0�hm���B�-����CV�5ؒ���i��|�m��3{%�#�|P~P�~Go�~DDD�γ>�]3��c�z�����Ei��i#��Iė�������/č9xO'�E2����ѝb��a.�X����/M��=�;�e%5(m,�r�T�Bڧ�����܍5:8��GGG��؁YX��w��v����H���
 q���:�^�)b���,z�n�}kԚZ�ۣ����*��*�����x��nǳd6�,SJF^�j̎c|k�*[�����������O��T�(&�w���2�``(��w"lhU�E��#�ڰ9�Gt�t��g��-f�����B�m�b���&[;�X�G��mm�3^�$49 ~��C^}2#�h�o~u����әw��D�h���� `�5���>��%����W�o��eG�� g߾}�1�꼍u�$FEeA-F��!���&��< ��XCBU#.>�Z��j������p.շ��� "��>�)&�ﻏ6b���-�W�А!j���<�z�4XKĘG��RY���p�t�JS�8g�Ϟ%�d\�
�l+*�?�L������jx՟�u3k���ׅ��L�bao7��AC�Ǘ����;,d򑉷�`��}�.����@a$�+�&�@i��k�4)6�x���6�]p��U� £s�4Ź_�+����BF��!��&`7b8%�^;� �Qi�y%%���P�h`	�Y~^�c����8q�=���|9eeD�
��+�::9�簾'����!�D��Oz���,%a�ElA���jq7�go�߈�;������
��Z�R'^�����W�^�D�`G���?�H�X�/�k���,T�'���F��R�P���0o3�ۦCW}�.~(e=��D��4}��y~ԩ�%9X�4wuy���*���K/8�k�S;�M��@4z�#~|f$� xZ�xN�-�F~�n�P�S���f�ʭ�K�_%�b�Y�ؘ�8�acc���"5x;�?i��DI�(�ߌ�,9O�)gp��Q�7ܦ��m������;b�o!!iK��m��f��8`�n4���97oy���[p�n�~�O��O�/��*��}T~����e����O��&��X	1��r�~��g*�]P'��4�Q�U�_���u�6�9������z���щV�h2�Y ��A�<��_����ׯ_��g?]�V��Nv�Kv[���D��S�=��ڭ�~��A��9o��=ū��/�����C�v:�$�V��n\�u_��3p��
F�#���;-����Qv}��2ڼ�ή�E������k+����?o@Y+�B{w�2Z��po�S_&�����s���މ����vq]]���E�z�,o��a���RDD�%싩P(�h�^��#�����~��&�^�vc��~�X$'$���������L��*���J�zw��L05X�qo�b����F@�����R2�m̽}kp�o}�h	Bϟ/5<T����_m2�Y���i�ƽ�fл�6��\>��4�Е$�V�t���}C@@Ӹ-�Xt��eB������t�������`�[�5������X�Z:��.�#Z!%��!*��j(e��_��s|�4E,���̓����u�X�������'�,��P`��G�5�q]��v�p���h��Pih'@�L)�UUU���
��1@g��zr�k�	cl���c�Pgp<�9$EK��89ݰ.� p�<�JnPpp82G&�^d.ɉ�uI;;7W�cU�L,�{T����^�-~X��vZ�;*�m�c`j���X������*@������d��~�,1��旃:��G��@kUiїaV��M��E�xڪ^.~�������zΰ@�?5-�~~؍�S5~/�r��N�6@�d%��@�cq�E6��h�9+��~
���2���៉B��1<�T�#괪*��5�U�99����~�hF�8��Eѥ�����eJ�����,Y��(��^�}� ��nb@ðid��,3k���|3��_*�덙>�n:ևz7�%������5��E��~bjj꧝�PL�i5ߛ^�����G4A���*�F�.AAA�:�]�~ �#��+IJJ�:�$���q��ˣ�v	�`[ۏ �.\�k����рF�v��p��߯�{���-y}�����atR�����#��W�5�l�w�#=O)H}2D��g�n���&]L,�0_��
/�NH�䐵��T2���<�}t��O]�����;Tl��{��1e��a�:�{&V��|E�Tn�� ���#����=X�8X���2-���Й�2���U�����J�l�7�������5����j\�Z9�%��Yf ��ZC�hML����iS3��'��)B.-�_�����r
ҍ�</~ �q��g����B$w���&�����S��"�҆��8����;���*�P`D�8\�뱵D5�<�]��U��,���???�W����$�w�y�l	P��ր�Ϯ)�)",��·ՇY"��#_<	s짠͕��@/g9H���4��M$�ώ���w*{��� �>�q۱E
����c�|9p�,˨G�3;D���sY��W:+�-����UZt���L#����׹D����Ÿ��~+�S�ɾ[�wuw̯��y(?�z�©`a��q���{��$���J�A���� z��(ʶ��çO�}7�,!�Aع�~%���D�6����oC�k�B�[�h�������|�j�#R�H�D�|��!���ˌ9��\t��ِ��p��=ܿdܰ��1�72��O����"W��)%��l�5�o4�����{�9��
�Xϰ���H����-�=}�w�}�ۗ/�y4$8o�t�٥H�:�vA��)B���޶{^�	���|�AW/nDr��mQK����i,� ��)�#��i�~��ut�7����G`%��+�ak�P��y��W/9洴�pP��h����t�7��3W����%�ħStU�թф�7���*�K�kM�kb}���\�E��!�(���� ���Y��U�(dS���Ä�UZ2�s��s����[�2PH��M�vK��JD��(��ɟ;��J�kW�C�~*���1ş��EP���-�X�Y�)�C(Q�*���S����jjhd���>�`_��4ڏr|��[�=�+f�� ��������||�p����6\�j���lؤ·}���_��U+��v�mX$f頓��t�K�/S���<A{�0N#����yt&�wA�рqcw誳���r7O�v/i*6 v%~Ԙr7���
l`.���eg'�'Y�w��T��@c�W�b]��|=�>���: +G�(�|�r�3d#Y,���7$|7QP�:�����To��Xnt���q1
���1�BN��:�4��c����N��c��!�N;1��+�kK�@S�x�	����1��C�{Q����х��TŬ�<����Dj;��0�`������	�>�l�>ɖE���ܾgn;����bȟ$��>@���_��h&��J/�k���ߩ����-�E�zaº~�)����1v^�Bå��ah.��u�J�
�������(6��ł�Oo���Qq�	l��[K}@睻p�Fu��e����'a�ӈ����x�'����q�r���E�8"l�z��GJ1w�?RQGw�*���!�ZVld>�2���ph�����W�sJD����� $��"J�JZ��$\�r��w�U�e�&+Z��~��O����'�s�� ���(O���..��VL�kih�IH2xo|ߛg����ai���=O�i���`Wd�/�ǆ�KD�lOߍ�8~�4���5��O(���~��&WʘC)�{B��v�a��'ڥ@;3�C�O��w�}L�;:9o��31⩶fA�!��Q
�2K�.|�B�2Ԋ� Iu�Q�w�b�3w(7��i��R�g��ְ4S_�ؘ�iQ�P��5r�Q�^Hqڷ�sfD[��v�G1��<����m5�Q4�$!h�rp��hTu��Ǌ����*�?��M��x~q��l�g�Ib�?Eبs{���{l���t���ԛFC�@�K~������`Iw�<=DZ��|�^�������0
�V����E\�jjj̖��7o�a�j,X!cjk�8���E1>PR���t�$Z���w�Ξ���	XO
W�C�����-���%��Wd����m�^����Uz�4�hE�̩I������f��j �B�딠�7��x���#m=�ͦ�k�����!�]
����	�u$og<��Żt����G��b�����'���T����|{�3�e5����B�T�e]�8v4[���~�����"k�Ey�v5��z�i�x9����zš�JG�Jp�V6h�Z.l�L�3-T%����@�طT�������$oW���>UŊ+��-�*����܂��h�͛T9Y�+��Y��t,ߙ�'������|uF��v�m������rB�@�ʊ��dfa���RQ�1��2��"�������g^` ,q��$�]���������eeT�Р�p-�5A�i4
5��e��Z��o�3�j�J'}� Lɲk$�>HQQ=�����+k2�����V�^���D~�f'�cf�H�[�N���m�y��L���j�ԻV�E�G2-nw�n�`M���M���E�d���
�(�dLц�'���J.���6t�^��c�VЩ�J��4y[A���6^������I��z�$�W���`(ȫJ�R��^���B���F��c�ys�o��Jg?F*��0��?�~��N��C����w���F���F�N�ɢUNsJ��7ђ��&'�_�v���dgԏ�7��f��O0��u/:Oayй�����G�Mv|w��Vl4y���]ZY3�`1����{���u�2�[C����t�����%���<�=�OD�0-���Z��n���&m�m��"y?�G��O�xގ��b�7z�S�k��'>����ȝ;SL]���n��t�����1�5������f�+�FX��^���q��ѧ�0A�q݁X��p���`���*ѬH%1��f���R��y@�a��ٗي��欟��o�x�&�Œ���k�iД���0�@�P)/�qt:�4��!��ɯ?����-g��!<�C��Ŭi�#}�3g�P�r����*{��%��1�9y#ݷ<�s���C:"��$��Iņ<s�DWZ�w�\6�7j�Q�E�&M�5\"_O��Ú�dC���_����:�܇�[+�S��]�Ll/�$��39njj�%�7}���K�Po��__�<��2���{���}X�+k���n���*Ņ�p7���bu��M�mV.��,����u/{�㥊�B�ѓ#2e�
Lp]�_�)��>�k�*��縇�8nc�<Ǥ�n7�>����H� 5��mf�f�]S���=�>dc�����Wm��
��#G�d��ͷ]�PM�i�3+�N�O��W��8�Ǟ�#���=�~O�[ߟ_�<j]�=�z�����-�Dad�VƊo�W�l^�g�?�ua/��(_�hƳ�Y��Wb�FNn,���m����Fj��0�x��虧/W�xļR�qC����h��������8l�8�T������c^%I��s��c������.��K�q���ϫ���+A>�="���$�%�r���]�1߲��)�L����1���ҭ�Q�y^(hb����r��q_�q�|J��b��W\{Q�(>~�"�:܇2�.y%l)��,*_�[	<��AH�����ҕh��������Xw�<Y\�KI��#���=�9��g�V�_�y	Z+��e������Lr�'G�Ep�y�-^F)֫]ۇ��jY���va�ha�8���5t�����94��.|Ѿjfa�nCl1��8T�6 ��P�L�k�:n˭PqL)ds�ՐT�0V�2t~Hǉ��0mwu�S^z�|wF+֢���K���3T�z�D�1�%;<���$��pM��D��(�UFX�-G{�b�V���%�7���j�bX0�`Qn�l@����i�24�(�*���W�|�A�b�v��˫v���������qNξ�P���Vt�������]km]�n��Q�bIM���s{Ɓ�CA�6��B�G��Ӑ�����Wi�N�q&'��S~�s�2��w6��3��N؝6�+Z�:���oc��E-��Z)���4�E@�
�0Vߪ�5�Z�-�S���
=x;l����K[ ^�r���{��.qD���D��k��X��uU�3�bH5A tޕ7�w��¦#pʫW-�7�h���L�=�w`E�^�b���md*r��l���\��ә�[�cm��ϴ;_���eR���B K�+������%�]��+Ҟ����(Ĥ����s� ϞIn���c�����1�
�acm���?n��o0b��<*�g�ض��'����XyV+e^��9�|G���x+,�nP�S9��+0��?��fߝ�Yy9�����^A��v���������,��_����X?5�� Otn���It�H`K��s��Z�Qd)�J�1l-�vy�d�
soi_d`(�մ���u32�<��_��n���'9Ēn���{L�&Y� � 6����4,)�4��۲6`LP P�%ߞ��ʦ���,��%���q��T���3���/1�3��g.�s���5N�9�Ű�?���v��L�H�6N�ϭ����@;􍋏��W���Ћ~�x(D=ո��.{d�z�tYL�rC���G&�j�,ug
�0��q�����
־�;��<#;�X�V�D[�[��[46o<94��Y4�f���l@�H;��p���nrd{�c���l		Ef�#Op�GVsD���.WE����.�t�������Q��S�-��|_It#RE�#�n��bI��6�|�Yv6r�&�O5�Rh�i3��c{=$o�t��r7��.�w������Y��D7��l���WZ��E�.��� u�{�]̿%��q5]�Џ1N��$+9�f��?|�Y�'7DN2�gK>kXX����2V�q��/:ܜv-h��Kg���H1<�>A��Õ�1R�O���˚`�Yk<ᝦ|��\z���LA��x?r"��T�7��y2s�У��T�h?��EW�[��/ghX��!�閌��5J"��A�!�$#]:�r�0R+�bٻEt-��p�59F�}�Ϗ��������cco>k��R<O(,�o���ˑ(�X����l��.��>r̻d�@��i[%����)f��s���m���^n��j1��u���B�9Z����5u}��^��@fG��'�_�:u(2<�_w����G|�р�Z���w�`�1�#��j��b���əZ��C��Ag��O& �����p<���D@7j�)Ж5�r>��wf�ʵ>%	�b�jz��y�>�7e�c�@V��!��y|Vw�$0?�b���-��=�mbp���+r&?&����D���ʿ�X_T�;�!݈͜�U^A[/�W�����,Y�k��=ٮҌ�IYwc�v(��a�\���+
hFTi�)�;a4�X����O�Q�����"��ET�2�%��d�a� ���֪����r=�N�_
�3�_>�F��Mq������wy�ҡ�'�dBIӆ\��U��
���?q���u�R�5i��x�"�V�H+�
p����/�5�G�x�[L8���W����混\ʖC*�3�(�*�C�ve2�������뻜��,�tJ�3kWG��m�"��!�K����Y��1���9qSU��L��-��Is�1�K��~��]��p�Q&a��gБ�~��w�����)���W�J@71�x;� �RK�{rXѣ/��."F"�V�����GZ6f}����qK�����o|�:��ϼ�X��-��WۂzpE�w(����Ɣ��V�I��J�v�cg�M�ݎ���_<�C ��N��|ϋW!�[+�_X�+�����$!P�Y��%Ӄ�m���@Qek9u�z8>�'=|�BVK�c`c��������T?S�b	�������J?���D��G�qBK�n��gm�v~�f�g	"OT���5��g���v����d�DWf�f��F��d��8�_��|�r��L�;�B⁝_�WB�{��R��9��3�����~���ׅ��ۍ��,�yϫ�֣8�e�Ѣ�|����]d�n���_J��Ed�/���2���(��7K��e�BQ�W�A+�K�(�b�n��G�Y��)����������6��|E��
m�����|BJ#�.Y�௜������:{2���u'����t����74|E�GBM��v�wS�,}��yS�����m���QF
*R-|�?�SكS��۫��AĬ�7�A��˝��$xٲp����X�0��6D��y&K;��T�p��:�r7h=)Tv�?^�%��3˷Ž
JK�	���E�;u4wK\��d|�B���|���$9�-��{��ذ�g����Wc�#�ԇ���\;��y6?	����h���>�c���#�OJ�C��|9��;_IV�l�m��ܟ��S<p�c�ںz���G�5��p��A+���Zp:��o/ߙ���e�H�Դԙ�����n)"�i咯J��D����)��~~�W����8��.Q����0�Eo�׏=et�κ���q,$+�)v����ce�J9��/5����V.�0����wqR��%}�[NHɲM�_˾/&�ޢ�L<�z���G&
��Sg~9���P��X�H�K����M�R�GЕ�{�[|,^�obi@J���]{��t.�h|;2��~�F�9tnsIRuk�w5�	"���c���K�Ƚ*��{�}���uRM��CcxB~&}mJ{֔��'pS�z�b���l�O�Xa�Z��vp�纻l��m;���K�R�֠�h�_Ϝ+1���W������-~G'V}��Y��b�~/1���,�Gv�f��5��$�{�ə^�s��5�µ�b��G��+��A����D�R�W����=���������ݵ=�;S�/K��DpmM���7^�:���{~J��9 ���O�4�*����W�\փ7����SӹR�Ɂ&XcP@���UW6�� q-z�#��=?0���[Ra&?s��3Ȋ�4�����X�G�$���>�"�;Z�����8�\�h,WGWؔ�$}��mΑиy� �P�5n��]#;�I�L٫��=Zym/yc���h�ъ����_��A��W��Yu��/�uÔB�ʷHgX}�kE����,��v�fk,m����UʡnB���֭�}�=b\g2���!Js+H�vL;¤O��ZK�-��_#��g�?�DڏPS��D��<�>f���g��K��K����%�&�܎������2cj[��F���mأ[ }̢�DE8�>��/��2����K�o��;5ȅ��-/���֞\Gx��P)i��;�;��Bm��#Oz��<_&�^:c��#$�N�KZ��T�u%�n��^7��4�[Ib/�0J�?lg���YY�?��un%Z�"zN�y�*���gBFGy �x�8���y(�c�ԭ{]������$Ez���,-��2uO����Ԗ����z������ͭ�2�|f.�!�0��C�-�ŭ�OՖy7���Y�m	�47���s��~KL7J�xJmw|\��N=�������(��}��P� σ7;�^43*�j�Z�EHфzDXj�����h�\� ����hH`d�"�L�}'GIS1�
��~��+U'<�vz���K��h��?Sp��O;ig�B�&{�e�z"%5����b,T�!eny�B��n'�F�x�*�Dq�����Y�E� f�6�õ9>7c��8�
�7�IODUu�����x�^,�I�N�T����Sa0��E̛&��˩!�0�'T"��/��|�����2m�?SJ�z��XL̵4b�޶ݡ0�Z?�m�;!c|��eW����&۸*�t�|oo���c� w}�~�8����<��b�Ei�C܄IO�Dߔ�_w3����<�}�~� �L��3�qY+���TP]*?a��~�>S�냳)�A;��$�^H�v��>/�ft�bU �-��iWٽu��* ~GjRs�X����Ğ`�Ocv&�F|�N픵��ut_Hq���7���7MFoG��#���7�=��)F�}r�s�3+������Q����qU՗(���V��Π�DS�V��
��w�ė2(KQ��BY�6�e@�z�h`ۖ�����q(}����� �r�އGQ9"�
�������0� "�C"�C�
JJ��P�=��HK�Н�~P����?��\Gq�yv�u��ޱ���@w�O�0��!e�դ�x)�� �%����~G�m+SֿcD�)ǒVZvԔ�*t����Ė��h��%�z�\�gp�α�������L?©�5}~��~����Ǟ�f�)�L03aݗ-�n�':��"�"$����n���U��:y�5\��a<ܳ&�y=���t�c�ܮ��KJ)B�
l}����ģ��k�D{{s�h�?>��ͧN�h����/e�0�t�Wa�󔨟���,�,LU��`���"5�Wq��m5��v�]���Kh���r%U3�Т��6ZQ���x5�Ek��Q�<3S�e�\�A<���n*3�	�t	�t${N^)Z����K9[髠[|���SeN��+�N9�&��f�Cts������O��;r���z��pFL'55GY_y|���������2%e��ק$��33Un<]n�	{"%�$�x䢭�x�sr����²(q䬯���F�ECfD�wh�W��F��e+��馧���mp4�~X���2(��;��n��'���?���y黓�{�����9*ˏ���D�DD�?��~=y���ۮ�R7N�|�#���_[g�˧�t�>�m$'�h�u�*G�F��tZ�!*a}�.����N��sŀgޣ��s_%}|�t�Xӿ�ݩ��Ԓ}���(��b�#���k�b-lY���j]���{-��iO�$���'6���-��������ȕ7k�9��ST�6o�#^}�67�֪��	�QU�JZKE�N^̃�X��앖י$a>P`ZXT�=��E�!$*
��"��u[okk{�
�����O��|�Z﹞t��d_�9���������ʗ�d�	d�� O�RSM���<Gax��X��l���� ������)6�?!�����h�η3;�͆�<�g��8V��qV�*��n���R�^����OO�~�N�G���4識�	�����]p@C�4��>W�`���;g;'>�ꙑ�J�!RIv�rJ_�5߇,^��-�KEdk�ol��Ő�_na7��2?�w��"��gG1%%%��8�F���S+���ȣ��67��糐,Yʆ偗����#��E۪�;�g�T�
���4t]�jڵU'�Q^�T:y�Ŏ<�nw�ל��k1��%�1GA�=s��r|}O?n��C�����������E:H��RƊ9�EO|=龿�;^�:�o3����xW�,�\wg����t*��cU�!����r�;ꍯM1L�йp�d�X��ϞV��v}p�������$��3.r�,&�h�숖�ꋲ-��7��z_m2�1�p�e]#�y��Žm��P���[�����ѿ����H�n�@���[����U̐٬��2����M����~��]g��L��z�;��c�xZ�|��Bx���{����m�$F8'��"�a/���no���ew���C�����@��aə�H�=�����{O�vT:�dcg�K�i�$��z��qKJu��Q���)�@b�С�T��B�p�h%v��:e^o�zΛ�J��ի�g������99�����i5�����g3126�x���{8_p��8�:LG�^:�ly��ezBpo����z��Tf�2_� �}�rm�D~̩nS.��㣍�X�C��P�1��-Z�n�g��v�x��:.�|�bΔS��fOr/���SU�q�	�癤�Aq��2��j;�w֣���6:kI�3��1�8����ڶ0(bQ��4?_�j������B�?�GG7�bg����pw�t^"nV�1Gm�v6����i��W-p�:����UG��l�߫x/XK%����|�;}��Ā��iB��FP
I%�J�j��K����o��HZ���9�N��s�MJ�oX�'��^N%��52����ٟ>]y��5��ٳg�deU���P�J��e*1�󽳝I� �����}%�膙z��N3nͩ�vF1k�YE1��dnH�e���R��T�z��~�؁�����VlG��D����:���X��[�x���tFW�L�s�q�b��MwC���܂$��c=����W��������xQMc=_mix�:+.-6�m�߽���|_�f�-�Vz)))��ϒ.s�ƨN�(?�f��$����l��G�s.���p*dp������߿:r)|���Q�]"(4WUQ!ϭ<�0"S��.de9�O��up��V�$i~�H��xW�QL�~7BG�Y/���Տ����j?z�X+F~�����+��\c�'A9�A-�����5��pB�^�3[��p!\��R0$�|VVpe��
���)*OM_i�2W����8�&$̬˲xn��z�j���q-&뤊㐰�.v��k݈����{̓���;�B���;�~f�U���.]�R������⒒k�q.�S	���XM��@C�]dӆSf�ˉ���Z	OxE2�ߗQԽ:���x6��5\z[h'�j4_b{�.
�O��ʦBBXs�:+��>g��V�Z�ІN���H����zO��E  �
W�"̨!�I[�g�;}��1���������&(6�����t����Ԫֱ6�����i�Si��L|��U�9�
�z�06x�����!�e-�������#�l7͠��5`'�\���5�{Xoc��;N���W�i�SSщ�5�#I�p�_�Dn]��''�=/}Æ'���Q���M�X����r��D M�q)��,���������$���h��̿��+)(���w;��I�5G>IUԷ�*hI�_�G�j�:��MR:NTy |���f{�q���M��WMM��[_����<�<łh��ݪ4Bn��e�u>����	.]xC##3vv����H];�#+���`AAI���@GG�x��C������V��s*UP�II���Ϧ�)�S��[��54"���B����з�" �@׬e#�z\���Cm�*��߼�E�
@�"����"5es�g�!�zg�ݴI��Qzy�L�rv��͛*e`�NN�5��t&5X�k��̏�/��(��#�a�T:�a��2F#��V'����}������ԉ~� �ڝV��\a�S�� ��7��4���֚�(}��e�g~�JKKsVB���F*J�5\\\
����r��[B�{i�h�GN{ss���`�^�����(��껲�&�q���Ї''0ؙ�i(������Z�,���	n���8�,�|�ljr�\J����6�(����lj'�<|v������8���g�1ek����w��^h;��?>�EşS��aa��H]'H����g�J
��mJ�|�F)x��\�\s�=�T��"��>&�yn��s�����^=*�?�IFKkonkˮ�#�l-�|	�ϢUt*S�ߴ�N��zff���`�i��Y�MLL�i�E�Z����1}oK8�>_�3�:��g-�o2���µ�YK��,@�m���U'��C!���Ly�X�)H*.�P:�^���X͛�����C��tez�� ���.S���F�Ħ7)-�Om`�,�iM�I�c��d�l/e�T��G���$֟�n��7o
a�ast��IϞ�e솲_Co�p��qy@�ϫ���� Mpʔ�٥[���Yw�@̇t~P�����4E*~�����N�/{�+9�))��};�P�`0�DK'.0ޕ�.���q��)ڙ��Sf?�>Xמ�t�̃Q��l��Š�)@���m��5����U��Q��L��?B�.��r��Ȥ�.��\�%[sNŭ���=J&���
*z.pgCqqqӃ�U*n��v	t���s|�3�ɝ�d?�'�蘘�eW�I鸭�A�.
���`�fS�����D(��Jj�yp��6�?"]�e+���p=	�X�'�ɰ�)�٩|e<+y+�5��l ���m�U��[i\��V�DIu{���b�'��J��m�5���T����Л�q����έ�������>�G����6���8�h��"X���gɠ�]�Q<�>��٫���[=��{x]�P9֊Q�n�'�D�`sX��]�#��OS�2� &���	]	;i+q�L�N�Y�0�I�-8s{�f%�;�l-�gt=4d��:�����n#␕=��L�S�-_��݋�}��Ĕ;0�=��jA�MN}C�9U�#�th�(cy0�$,�}���eK`aӅdq ���d�B����_K��k;B�ef�+74)g=�S�H0W^�)����PϠs���,��W�AF�;f?{���2J@���r��{���g���od������ȶ����Bw�N��u��-��<���X6NH:�Ƣu����㊓*�cI,�I��F$+�_���L]�vH��˚w������R�G�JO��(�D;G' ���B�#t+L����ǏD$$��6_@�X;G���ܬ�CQ�y��F)���<���L��6g�1ܘ]-��&�_��`,�z�;V3\�Np]*� l|����I	 7M*2==�e.9���T�],����`�u=������D�=��w���:���R���u�Jlly�E>h?��&��o����y'�����X�Q^��7�v�^rY����xql�k���� ���QRA!�>�!�4�=�!(

��B�$+�סZR����e�*�k�
�������y[[����@�dC �2~�h_����	����e�&��P.l�h^ņ@���ii�j9���/Y�v��a�L@�2�����g-∁
	A��~�e������Nl>r{��)4bU<����Y���-͈&��a����#��]'�PS4�j�f�o�U�>��o��e�ͩ|5"!a��8���w��SOp�Ƃu߆BhF.��~��G���;Tj�������OxC��I~^^Hh�q��h>�V��ݦ��ϣ�Q�۷Š��s����G�gA(�L9���}��0e>�t� J�W<�TW���f���������@)�#��à��#�TPQ	i�����k���4���$��c�<��y�����H�e�QU;7����{����4h&��8�o���������z$0��F���~,�3�|>Z�?�c�w��Mff�s��uҺ�(\\�|0�$���X�X4]
������'�.�N뾡hYw�ﰥ����wƵBJv�����%^{i��O�����D���;�?~�o�v�A�J�a���m[�0�����n�.w��>�<��./����Yٗ�5�ώ��*֒��	U�xEH�t<�oM�[E����eF̹��
�M:m�$�nR3g��������9ם�O2�v�@��I�y���l�_��'#�A��&��A9j>E˺��K#�aoߺ7C5ej�;��?��V�4:������o�Q��"z�||@�� �`&��:�����	a�}��B<p�^������N��ged�EEEe����8w&<�O7��f;b���� %]Lc���puv�m�uo�(P�#�디�������c��^t��ӭ\Og:ߗ�WP8<UhgkUs�\�9�(D����/pT�����歳���Z��rX�����Ǩ�E~�����Jy���n�e�6�9���,x>V�$������/ĭ.��(_��X��%��p�[m�.�U�����c���ɐ^EFj�H�9�,�������//���:��(�0i%%%R჎���V%/l])�]�»ahr�f��f�z���A����2s �333+��������4⺜�(� � %������0l����C��T�n�Ny���0=��(�vg.���j/n����z�g�O�r��JHH�W�k�҅��bE+BG^
�ꯡn)R�6�O`���J*�:	�l�C)� ���>�~Ip�x�oݥ��f*�����N_�#������UH����d+]69b�7{�;�\����i�����B��j� ��I��K]3-��_���a�m="н��XHt����٫�9(��y�c"��r����P�'vQ���O�7�g~c��:W� ���Q��&�<�lh���3��@�#cG������O]�<,ii+|�������ի�1.w\�n�"(��ǹ%��ޝ
�]�^=�� ��͆�H8;;;�� P3��E�����Rn�̠5�;&���'�_�*:�}���~��Ya𘘒2�>F�?zA�x������(Y7\��}A kX��Y$4����3va��P��3�����D?ck�>_������, �O���������l&���lb�����6�	��?���'$$t�z��7��B�I�7����?g�`�v��ω���'���+�ڿL�O��w<z��UlUu�����&�ݻ ��!uEP��!�����"���KG��	@AG��v���!��v`�@W�����K ��=555��V��z}7��p�&�����ng���;�2�IL�խ��6٩�t�?�"6��>�e�)�\���kޯ�W��'����^I��~��Z%m�L,�5K3������W���x���Gh`7 �e �)��莾2#Ϊcp���fLh(�	+����d�p����֜��H%�N�y1@i��OC���\����{(d?����o߾�Jw\�p���`bb�����+J�?~�C�5E&^��]P��0�Gy-NDU:�g���ݲ�
����U�T$%�]fվ�������2�R���D��ds��e���A��o?�@��C������Sh��Flq�;���Y*��ۂ���VW� �I����4cFc�{��A��ցG��_�N4L�:��àZ�ȏ���Y�'r�h����\s4�V��?O���J�ҧ���> B*��c�A{O��H�Ha�*��T� +A��ai��(҇q2�͛�j"���|�N�2v��Ȩo�
4N��v�0��}�t��v���<M��o��u�_��G�c܎0�-�2C�Wy�gf����C?e��)gBȞ���峀ׅ&���E�9n@s�|]|λ�A��Y+��޽���-Y��+�������R�Ӝ�Ν��
�Ќ��؁��1{xV��!Tn/>�w��ֆ�
x���E��ԗM�m*�?�0n[
�2ƕ����H�D��Ѥd�9���c�h�Z/Vd+kQK]���L.��5�P��}�9pô�.�I��N��{�bon/��K���R�(fm����en5��!M���Y��$���PE�]�!�}�����:g2�455��@:�A��~�>H}Wl��T���ru�������B�	�`��:V��G|jS��c�@s=0�mk�q��2����Vk-bz}�0�o��$pQ�æe�+d.0/��w�Jcݓ$�嵜;!�ԙ]v��PQ��,�p�A�"��%iY��ǼO���:ϫ���?�o���?�N�Z����AiD:�cR�?}��9�������	�)d<6�4b6	��`��);۱A�>�^�ΔT_o�/PE����Ў�,%�g��N;�_�-<���k�(=g��4�Y�*Ğ?��͛N�ԄQ��{��/�J�&���ګ�?�F��-Gӿ�W�ɮ�ʟ�t�`m@����F�������2�33�����-��Ш(s8t��Kr�0�袬Ũ�H38��FZ; �Ƞ �	#�"S`8�w{�Z��s_$���`�J��)����G�Y������^a��S���RJJj����-'�δ��I�����3��MEG_��(wX̨���u�ɝ�1��(S����|�fN
�����MvҊ	�گ���58�i�<l���>�����i�9��/ t���c��|�r�s��K�!��d|jk�_� �g9��.����:;`N�TGc>�2��aa�	�ouuP`J��e�L��O�s������ϼ�g�8�v���.Jq��w�u���#��I����󞧷����Yj7C%�&y�I@�XRRו,��o�,UE�7�����޽{?]U���S�y�ڀv�_�D���c}���YYFF)�l�������y��h�k�N+�k��U��,���Z��Q����J�����+˥'a^����#%�v�Z0��B�.��B��1��3� (��ǁlLL]�g�i9�d@�����:��2��׀���X�q���M�$s�7���nb��T�%e�Mt`�d�9|0���8��<�hg��o6U��3wbJ_#B ~�Lo��a�1L�Z��B�_�f�&�G�4VH������[��������x�v�ܷ4b���9c �̫�o���՜c�\�ǹ���� UJV6k�z*ݝ;P}� �k�Sd{�$H)()��h<S'��0�m��N^T1��2M�}���cL�n�U̜��'I0 �CK�s�y�$�
~���t[V�}��"q�g`��(�щ�V��������%�t�C���B^���{#|w�e���p�M\/*l����)���£�1Vesw���`MH$5Km�M���y�.!�͞�7�0h	��ߺ����W�L�r���s�n�J������˓q�++�ec��R�vXǈ�?_��V*Э/��h���k������j2��=�Q�툶���B�O������m��^��k-y|1,�-E�QӼ��n�"�ksp�l%v�5q�Ń?[�T			PY[T3K�N�R������M2���-��>����l�K]	�UK�@e�(+>^dnn.e��Y�gI��^'0�J<ʬ�3�oM-2 0g���}������m;��)k�h���i�[�k�������kx�Mb��с�����d#�^3�6ו5T��=��H��5
�b5��+�{��;}�˯��֋���S�(����1Y?��UTټ�R�I�D�YX��0<q�q�\�n�|eS�Y��M?��^��0=<�E�,H4�bI��Yu�v���YF��(��r��o�/�(�Y:�=.�+d\�(Զ��.��X��C��^��Ք�>�9h�2ٮk���ߖa[�W�U�+��Qop��U�VT-s�2e��B�r�՜�=���&������n�O�Q{l��r��c+W��e�D.���z#�Z e�܈<D�
��J��2�A˾����-dgX�Un�:�3.��ܮ�t��!X�&�$>��<2b>��'`���ޘ�^r��$��+	Ə���ѣ���i4�,x�8%�))�1���n���P��G�?r�^�V�A_�iǂ���;�5�%lv����R���i��A�L���vV����xI��{��ݻ����-�5o|% e�Us�E'��>h�3�<���k�������w���|vnm�<QPN�B@Z�0y�?�
������5_��G/�t�@�DBe���0�{�q��M��xh1���9U$����6Oq]*mXUlH��i�}�a&;�@��#&o�8ם:o��w<��я߬��U�y�6UZ���=t��+����g�l[����I�2��u��3��}M��T��*�g�[�*�RD��i��V%cg�R-��/��z�QY���wA��}���Ơeh���5>%�E1��3m1R��h�> X��q�EP*d�V �!�n(�;�[���˗��8&;��^t��;�NP�)�� @4����񵚝�~��2
@���DF
��[��aa�tڛ�����T�<e?���\�)�ں"�&~��T�faׇ�bP�%&!��e;���B�;��A�YP�N`?B3��C��M��9T�����9X��
���hTSQ	�8PI���;О1�������m���@�4дR22*��/�z� �7��>�:�B�6���3qK��wZ�\��R,U��ٗkjB;�*����ʵ��j���
L�d�,xL/�SYo�o���E���^$���M��RoL��!o�R�6"̫_�>Ѹ����R���9��wo�v�0r�����(D"ev֤ФST��~���6t�locζ4Áy<Z*�b��J����Y��hO�he�A�29�22=��
�B#��CJ{8�\�l��p��T9}f�p�ט�Sx��;72�>��i�|��l`��鿦�����%��aHT:o(���Bu��kNe�cY19�22-9��{1�>�p�'t�ǘѪ7?/4:~�Lù���jO�Y�u� >��4A�p^���;:H�U,0鼥�4�*`���t)�P5�a�(s�b��YfT��P��٤�=績LN��25]G*�G�S�b2F؎�0*����_,���v�r|�����L��] ;,�D�<��/�y��k�9�
��q��/�9�\��=	b� ���K�Y�E��04Bn�kx���?F���O(,]p=��ۇ��.N�6
�*.2Q9��ʑ��T �A�.�p������=���U�g�� �P���k���C �鹹�O�c��	Pt�v^���NVU݁��f_c0=�����!L�)ɦ �4��	iU �&"�;��J@q&Lmu������R;�[K��(���S���`d��
 �z������a|��}��M�Ѝr9dԮ�E7&�r�#oc�bX���fYW�>�RE��x{cg"p.D�^DM��qM��E _�XF��["8Q��=&1MN����� @����o�/��A��=\��@� ;�K5�o�L��E_rTL*�#�o��T�*�q�[�`0�P:h�\��`�*�1;��j�Wm�����U(6@e�U�0��ZOmfDf��fgg������#�z/��c�V�].��	�҄	��h��lS]؄�b,�����9y�*����3�/%Ezf�h& 4�|���+�<�v��_K��� .'��v(�2�"2���eR@Ũ Ce��14�͢[���;]9գ0;'xho������:��������x(�4fUn���j����-Sggg(9T:Iի
�QeLmm-5��\p�����d�� M{���	b>��]�9��<Pu �T��ǥ�c��@Ȟ��A l��$��1Pq�M`|�I�����L�R�����к���F�U��Gt
*��:��Uĭ=�hk[J)+:�W���Ⴌ��v���#��f:���a�m��ƒ��.W��~�h8��j��%��y�J��[�P�\(k�p���]����K�h}�fC��2&e��QK��m
��A>Z��k^�`�M����C�'��Z�^�>BM[ۼ2����4�4q��О҂CyMM�������[�/3ݾ-Dx��'�a<P>r(��?~\s�P	(��B�CCCT˝�v���κi�$��F1ݙl�?��秪����"ch``$^�ZB`��
j��� #77`�Νn�4����~�?_��v����̵��� �==N�>��ֆ���&~Qߠ��`����+n�����"�W�� ���r��5*�eZkL�C��!�â0y��.�d|���h��R��Y�_������� �Q�V��J�qE�������Y�*��"��s�C'���~��U�H�C��*�W� n]eu�ǥ���hXI/(P� �}|n��dK_�r���u�sۋ�8��]�z��NE`#ж��L��j��������2���<=!65|��y��wd��PH�8<Tx	�څ�{���'x�6����}��!�×P^�tT�w��M��Ha�%+�פT?��搛i��6��7��_�1`0�j��x�����6_jλ�>?�#��k�(�/3��]��{���FO�Ӫ>Y��<��vc}G6l�G��0�J-#s���X��w��?�}�\C��iK��\L�Er���i�%e�>ǐ�2ұo0��_�S�̞t`��gA�J��H%n�E�TЁS�N4T�*��a�@�k Q�o��N��11��Y��񖆖�k�����AfS��iN󤜙!�xU��_�a^fІBf{(�x���F��5�����X�ɦ���x�u�E�69�&�KF�[���y�9]JS�u���1~r��1Ẇ,�v�I_n�jg�O?2~-��;�5���}����U�>i
�6�պb���D�;�z�UA�˹�sf��I���?&Z,�6����y�b�3?��[�~ H>yu�;�MI����y�(�}��Q�k����)�NI@���4�,��г�������<��s�I��p�x��ICp���>��������A��ar��c��C"�0FgA�ѕ�D=�*�/��H��>R-XL^;?���8�[q�'��R��~N��~$j��9�_6o��<�"���a+5V.���-?IB��_Ŵ��"z�=������t<��Ϙ����N]��(��V ok�/ū�"B�&����Z?�m��g�jJ ?��ǽ'@q�<��Hc�3��m+���y��fL�C[��rx�T�yʚ%z#Sz��3����1�^fp�o�=p(\xӐ@��G�Y�$n�!��`��9CF�u���~]* $mHtt�y�5���e���h1�f�\��l�8�v��ȹ����S��Y�p�}��KT��I��qDk��D�m4?bjا�<_��������ע�Q_G4Z��Q���s�[I��S|m嚆�>��w���Nk�J�[kf�]��D��PѸV߯��IL��P��D���QjҜ��z.�Vh��UuY�'��TB�hR;�ghC��E�젇dǻO W�Oga�z��F��lV(��c4DZnqM�:��oXD�~�ǒ��+��Ъ����y��*�W���GU��mu!Ӣ��]1�/���|�f��b���w�Y:qx7�+�NR����{
���LU�QZPO���f7���^	�y<[+O�b����zy7�z�|1�U6�bE'�G֜_V�/>r�����m��y�y���qc����L7�� ���j1T?���]�{�ȯޢ�1J�1W�� v�a^u2�^�Z�%}��k̖i:_��}ON<|���B�Z������8��z���c�:GQ�]�e�Nt���O:�
�Zk5�T���_�{�u����[��\�IةG?�b�4�	��δ082X��Թq�zn� �t�����^�ӂ]ب����=<��꣮��sng�|�(�D�'�Tb� QT�ۿ����\E}�U��S���,�� ������3=L$XP�<����'_����RĨ�t�Ǯ��*>��T���|]�[@��Bh���c_A>D}��]	�ˡ;�:D|a�(r��������|�G�A�h ������\*Z6�ˊfLJ�1�I$Uл�����+#]Ӡ��EK���'j$Ga0�7�Ȝ���+ оta8��l�fP��%�$�˃�ٳ�����zk��?gV��Q�zN��R�|x{�GS�)]J����@����[QI_���z�?���e�H�>7���!��k��(0�Bz�'��?-���/?,>[ܣP�>5�~楿��J }��-!,~�oϓ���NI�r��O}Y���aS���Yk�?m���O]0���g�����Z�&>`\�e4��C����W��~��<�w@���T��z�$y�G�⨵p�̀gj<��ǻ�B�l�Wg��5��&b03��jk��i���#��	>VS�'� �go����&vb�m�Wy� �C������WF���ܯ�h���QN�7����2�%�l���hМ&Q�,R�b���z��v�OL�G�vJE{O9�2&ND��j�"r3����~>��H���^{7�j���^���Pw����:HBП ����������8�`t�vA���/�Gw�B80#\�B�^p�3;u�[�ߨ͠#0�~H���z�Y�B��*l��h���$��Z'vdr�9NA��#�z��\q�$����a�p-��u�G:$���F�)���[�,�0��h�ӄ����ux%�+���w�k�A�OSXh`;�eq|��/���c#q�������W�g�d�S;���3��i8�.��n��jY�}b�)B�b��Ӿ�U����ζ�"��4�7�_�eIO+���E|
<d����לG�EO��5�#�����ݖ�^p�}e@��Qc�
>�;q������ω�tI����D��xi|�Wʀ`D�ԎA:���?F�fi�|d�}O�&4}�<u5�ͯ���� �S@m�R�Z������K�_~ =�(���4�J&x�1�Cs���"O�n޼s��HPr���1��p:��t��6/8k��b��/9~�l:�D���k؋;��7FPK�#��wB�T�p�3�nn����`��%�e�sLa'�8�Ϝ�`�+��b�r���4�A�If������[���,B������ݡh�է*£���ܦ��ϖӕ�����>;�u&=��ԙ����D%���M�v���o���G������_8҅��y&�}����-/���؇�O��MZ�F?�dk-;c
�_��.S{�|���=?�
5�Dǫ���u|v����v��(ce���p���0�/��a?JL�����J�6e,�<f��Ӛ�nT�O�x�{5�6~.-����o��d���B����4=(w7ۍb�-
�*E?�Y��|O0���V�+t���*1!��]�O
]�ʈދ�)��aޙ�V�]Jo��z�����75_���l��}�3�N�D"�Wv>_��0&�B�P6�g�����<90$�%�2D�R
�5!/p�H^
�3����|�S�����3����LMer�	�q�k�_�]Q~�2۩1�����k�9�g00��eb�g��l+ѧX��_�MBmt�AT�힏G�.�K����?V�n9>:3s���^cV.�禾8�w���>:zo��#�i�����0�3����_��H���U�t�9�����['>G�\���Ύ����K�{鳋x��.[�GnܦV��ic7�Q����3h�+oB�H��t |�m	>%j<�v�k�ve���x�[�������|ܲ�n}��-��5#U�~�K5C!��9�ش9����;�y�=z����L�u좍SAQ�--�EA�Q���0�J�?n�u��9��Ao`t4=�3%�q�8�%j�@�x$�*�g]i-ͭxZ��������pƩ����������"�݌���&5Ra�dN�[B����Fu�I�o��]R���VfX,̸z�Oji��oڭ�h�-r��|��"�s�����}�E����B��~4��3EcϽ�s_��\���{
ҚB�W�D����ϴ
�/
y2x�IΧG�K��j�3��Jta�Q�^M3�6�u���q�("��P�n�����-M5�%�6�˷�&?韙�ĽҞ�|�;��ׯ�5T����2�u�P��ݷ��Ԯ=�t[����X��V��_o�� _.ճI_w�^��Y=M�PU�e��������QHu�Px�>BQ-t0�"�����9rYZw�4��oThWI��ʼO�Bg~9O�77��n8暵~>_��L���nf}��SQ���^UXK�z��κ������{�dɦ�;Qj�	��m�F�C{U�~J�/m������IEtl���3����6�k�/7(�����Q-q�i���TZW+e��"Km|�]�΅�窅[�߭�c�x����=ףlvn�Ĝ��+=rc]�Lea���6F�g"'���/���
U�o�V���ی�g��z8�RN�v�`*�A.�,��j[L^�͔Xg_''L��xmv�i;Ayb�α��CѦ���q�[
&�żQ���8n�pt/��[��o���I�؁������w�����/���Q���1e�]=z��D��:�#������5��j���~\W<j#"���4!�_$�����[B?�{�c����'�y�V�<h�µ?Ͻ�����Ҽ�	���G�<�;r�q��7��������y/�<�>+�wm�R�-��F{<��u���$ò�e(���Vvu��� �v>�z��Οq��� �}빷�	$��DsR]�5�kb�y ���w��$w���,\]�d���ov�e;a7I%n�,�����2�Eƴ��x���	J.Ҏ 7�Rv&e�	��V�����G�S�ۺ�j�� !��,�xg�?�� �<1�����FFTM���褍�h���?|�����a��.�%�ݕ�F�M�\�R�c��h�����}1v��͌v%{��9n�E�!�͑���F1O�b=�_�E���˻݂^mb���߭psY-�%�pVAF�n�}վ?t���кGuv����9n�gr��e���<�Ke�M�g�(�<o�uվ�e�d1�FU�F�w�+���#k��#�cx�c�O�vo�ޯg����w �R�FD+~��/��{�	4�Kr��:�=��8�Y�s�gB��5�3��EO�Uj�},o^:c�{����N�$���k~&����xDA�'�Fn����M��S#�����Ky�#��V?N�+�B[Ԏ����"rt�`ZB׶�Ү<H4*�!���.�p�i��V.��l����T��g:48�~�2d�K��%o8�2���;qDe�ly��3������g�6�����JK�2w;7�D2P��Z��c����v��w�����D#���8�`=y@7�66�8��5$HN��!rA������]�`�`�%���73| �*n���@Ӭˤ��Ye��.7��?����h�1�����`�>�h��ے�Ͻ��K>K�<#�=N�C���O�a�J��[&f��(��,�ן*���2ɚp%I��1n�P{��6�U7;��R��.�}���d�?��7~�x�#P8�q�м`goY��~g��y�(��.���:�k�d�%���:X� �7�t�ZO&�)�'��/׽8r�8��t���6G�7�`���Xx�}NQ�,;X��!���lg���8�������٣����������S��4[��Qr��nK}��_3ދ��t�P���y���RΣ�#hr"8���]�������wul�>�4�f��.y�X��} ��{XRY��+�\�g�RY�Ԗ�a���Vr���	0<_W�]�ʒO��`ҩp��{�l��z�����llP��SR
���$�S?��W�w�����_��k�f���������Y��FܳepZ��AK�B}�5��t�YCN��%+�ym0�wq�m�*rnntWXXNrV�r�y���gI.nK)�U���d�,��
+m�z��=�GYH.	w��,X�S��$H3}�i݊�l���a
������Yƀ� {_�j�I���&��X�Y��x�����C��t�
)e�sc������խ��O�i<���	2���B��}��;7{�Q�6����v��څ��X��p�O��eGK�8R�<@��ѕXҙ�x�\�5���F��M}z�hƊ��-Yy�;=��TT<b���ե����j+��w\Qb� ̪� �=�7�w��6O}��G�]�3��}`a��$��`���,.tz������jֹ9߃zʼ6�ny��-���(ZSÅ��|��t��Ҧ#]����u{��l��5R#��7�3�7_���֭G<������Q9�n�-�V�b��)6�(҆��E|�|�^����붠rO���D櫻��7T*di:��M����,�����ſ��z�
(�x�AcK櫢�	��屟n~S>�j�7����cO�s㴶 ����Hi���v4O�;����[Y��`�f�-���6v��mvqjЇ�]��N�P�
� Ɵъҡ.�ع�d�dS8�'�g�#n��ir���h"�c�Y訲z�O�崁�ŀ���x�B]�������8\Y�"�:n[aa�mr�·���2~M��z(��ad�-���Ɠ��K��>2���������@Muk�Q���"M@DD���H��.�D���+��ދT� �t��Ѓ 5t����+��L�q���Ե����Dq���w�����f�͗���ML�L���� �b6_�}r)��ܼ�$i���Z�`{�&�>�2���V6��a*1mX�������-��V����}}9Rk�c ���~�M&���>@D`^�����S% _�����۾D�@g˿���6��`��o�^nn��m�<,Z��֧�fl�Qyfl���_+ALfj�6AɾP��-@� %�Vv�r�jv�]�0����Oh;~2�w�K�������uT�Y��6��}��qz�3X"
̼�_��+������<��k)�.׍�[߉��31�49[x-�����z@��%Ǜ3O,����>���c����n̾�)�e9R����l���1�"��u��ý ����,}����8������~��~dyv�ϢH���0�i@z/.0\��`/�t��WK�/�ڃFSd]� ��=?/��j��)'�J"������|4�1G N�1�8sȎd�������0����֤Sf[������,�bF>P�Q�m�t���E�_���1M��"@N权7�S��SR��Wm�ͭ����¯E�*����6;!a�w �����RF�Vğ]Za�
�&Eb]�Xaez��P��h����b�f���Y�����\y!���RU����R���D��n��d�OI�4��ծ�5ԍL���O7��8��nVy�=TI.�������O������)$����>	bylK�`}b�ȶ1k�#Y����	�>�Gg�n)���
���[?B�d��9������DgZ���D��?X(3�j����8��D��r���ݯ���LrpxU����!q��	b7�?��]jϠ]��V����E��G�~����˲D��JA��O����8��4GJx�_��V1F���[f��A���k[F� 	�G_4�S�--�.���+O����ٴ�S~g�%�Cς����@�����Y�����M�1�%F3���M<��W+DP%Z�����m���G"
&Dg��E��"���<��/˄sI�w�<�Iv!�?8���Oc�r5p$P9�겙�u(Тq�P��\N_���cd_p��:��:ъ�ݳ��;�r����8�s�Z�����R0�۝(W�������%k#������x�Ji}������Yb�x�+����3门5���o�j5���{�F�ub���A��V(����g���T��yfq����tt��^�A��#l����~�����z���Ϭ9	�n��
�"t���Qx�{ߣ����l��m��H=�w�#9z�����C�wD�)�|����ʼ�;��_�����1���Y��I�m�9$��|뾓׮olp����f��X �@r6�nI>w��¥*9o2�|����SN���jE���n�c-t�gX� ��F�l�1�o�i��6�u��6�m*�.��� ��"���ٹm������g���෈�<�k�ȝ7��P���Nz^�2�0(Ϙ�z�/�����ḅ�#pbӺ����/Ï�h$��>Nu�O��*���d��K�$�uüp��S�3;gm�-5S%��{;��G��䊱q�,%ƺQ,l�^��ϙ��\�f�~����e�q&����j{������zM](*�!AD��k�@e]����]�Ѿ�׶��?�ߘp�9#[�C�]��.-iSd��}�T�s���9���o�fFeD��Z�V	������oǕQڙ=����q�o�����<�	1ŐI�d/�VP��jS�Wո�r�F%l��z��/�%,�w�c�Ր�N��ON�pO���>���t5I�ɵ� 6�W�J`��6��]I���3�5�����-�צ�XA����2���?H§�����?r�]���j�@皘/��F��9]�]/�)c��'E�e޳,�\��`! ��J��x���ڸO���N_]��W=�8�S�.
�BT�\����<�������W�d�^~녺ףGWՔ1�w!n��$�aP��'yT���;$l��)g+mF����;sy�Dl���r�o*���uA�;ux��(�w���A�����"@a���	0ϭ������ ��e������g4�L� sTR�A|�	P�V�J[bzL����{�5+LzF�~�]�!�<N�I4T�'��l_v��	�;w�����%J}͌O�tܦ��w �� ?��+9gEe�@�A#wq���3�%
 zG�0C:���L�ē�|��+'Zl�KEتMV'��B����1Q�?P̯=�^�R<��V�>	��	��\��ܿ��8���"�vy���� ��Xw�#FT�J�?Ȅk߁55�J���r6h��Ђ��<��_�L_M��Q7Q���]�4��I]����6G
��!�%�N�0�ĩ�|��.����3��E�e
�`�R��31?��P0� �mAP�t��	+oA���I�mQJ&�����^uf�Y<����C�.. ,GW,Ӷ���-a���?��n�Q��]�buS��c��\�N]���1��0-����}�-gD]��4^��=�BV�uR�C��u��'؜\��z��YC�F~�K
0�d���X�6�67-��D9v�`8�<�k�KF�Z�{�7H1��k��ű�#�Ό=.�.!�$L�����'�:����ME�Q����ɲ�낕"���/��FD���.�(�1�V/1PFU�ץ��z��'�2(�`��MY㎝WG�OO�ț�1%��V�*�
��;V������fA�TP�$ى6ޙf ��`5ۄ��(��k�җ�9:� �/M���:=?J���ʵ!���B.�S��b/��f8� S؏Dw�pIW���?���7�sf"ց�`��`�\~����?c�ھ�Z�� ��P�r[Ɠ0G��M/�|��.�LY����=r��~���B�jN��*��A1RDN���*!h��&�`U�w�Km��& �&����1�D�+�V��/�X��NLg�r��֮�����Փ�͘���.
#����w`(� !�#��h)!�u>��&%�CZ'�<�Zk �Kr���It���C��h���N����eމl�&¡7�)V�n2�\D x7�41�`� �
MӀ����T��q�m��Aݐ��g`P��l�˺���}u�������U��'je�/L�]�p#I��͛el�=��hB4eY��[Vji��7�(S�%Ǻ�y!��U��,&�ƚ��|��@����[�������	���E�G��!Y�唇@��|T�>@k�L�z}3����aT�F���$��!�DP3���<q�^���.�oߕ�١��%w2�����z]*��3^��jw͞��2����=��N���h}X� ^�T�_��Yk�<��V~�bt=B����G����.a�Q���a�nģ��IH�.K��w�Y���s����E;�MEO�x���M��e[�R�>wc7��� g��&�����$8&*h,��ZoՎn".���m>�v�����Ug0��VK�nd�A��B��onv����-��sL�y�����η�
$C���C)F��W6�֕^����㱪�x�`�@F�m1���c��V6Ѭ�6||�}ϱ�K[Q�Ǿ�7����G�A{'��ktCf��{��� %���גվ��6�/H«P�3�����f�������79�@D��A̯*�_����ei`~c+���9���}�_2��u���˯~�IdÀj��טq���Z7����r=�[O���@Vht�u����&�8,���ϻ����C�m��Q_����0�3e��ru���+�~��P	y���E�i����l?�.�+e��g�Pa��v��j����2�Z�>`ҽa�hFJ�U�=��vР��K`�1I�48���8��v[ru�хL]�>�/��I�c9Z�`>r�j� �re������!��~��Є�09@��uC�a h��r�3�MgC�P0rE�r�H3t�ָEVT�vP���;fB�������Y����{|��z�u溪MHK費q�d�p.i������ʥ`��q1?b�*<��Z��o�����z��M��A�2uaJ�O�;�==�*�'��Ӭ��5��aKKߥ�ї����S�c�5.�����Փ��a��F���Ȭ΀R�����<ն��
�1BXHCH!
�9_�s ���sJJ}�O���JD��]���h2�9<s�J x����#2*�YD�2r�W塡t�VS�bba��DN�tsJ���ص���R�Ŀ���C�2�r�P`�I����AeE3��`�M��S��ԧ*�����z�D ��MJ�|�E<I"�i0A++r�I>nb�W`��;tA�L��u|���]��͡�⤝aȟv>�Ēg���S~��v�&�'���}r�n鏌�R����-��\�xRmh�����)��_����56G�L�-�7vح��C:���Lr`��K�J��5����OV��v���C�δ�f�3ej�������}b��3A����`ѩwŐ���R���T�S�6��MzԪ��Bb�va���%_�h����8B����ʤ�%v��)jhZ�������bb�zU<����P��0�]֎i��ee��+�y�c�un(ĸop�6�����:|�fw�'M�@}Vhܡ�Ս��a5�vW����M�%�{�=�%�������k��c�����|�W�p�����<U�����!ccf@�=i�Ӓ-!�;�?)z���[��V�?�G^����3���^�e�U��ۀ�B�0���U4j��j��^�0�5E�_�z���G�{����Ժ#K�tj� ���֑�.��c*qP���9��È���=+�:9�D �ȴ9_�ȴ�j(�����nMvhY�FN�V�6�/��sy��~3O_-�_�ڛqΘ]Z
AL�pwv��s���+�`�C �r��G�^��׍	�l��('կ�\6s��F�vj'��,�4�jT0��$\���b'�묖ҷ��?���m@/z}I�Fi4E�,G��V�.0$��C����ϛ0u�����6r�n�6Os��/U��"~x�ă��������Vp���MI���,\��Y&��:�&��C=�K����^ӧ�����@��+�4q�&����t����\ \��+Z�У�w��*�.��g����>�5m�N��k!b�o��:aM��lc��$@*����y��C��3��$���㜍���Vٞ��m���W�z�p���K�LV��s�{��'�&V�=� 6J���Jh��g(��/Y�"���	���N.��%Ѹ�
���m�`J��-\�<�`t�i���m�'�����'/�Yg���MȾʆ�פ�l�����Ax����b�X$|ʩ����d~0�Q��H]��j�i� af�"��ѹ�n�h���ݬ�M�A�w�&�C6.�4].ГX�5�ĥ�z�$�S�)��6�0�+A��O�Ϊz�c�j¥�Ϧ)�z�3���
�4�`t�r��7���SH��0����zD��V�2�����=��˥���]�R`ͱ�O���[�%�-5�E�{}%�Rð0����V`uB�z_nO��\��۷�Ć��>�"7[��;ۯ�K�{@\s���}w��7��w�y�k��O��/+b�s�W6���':����cx'z�)>�}�jpֳ-�%�Y^�`0�Q��<�@ �iZF��'sD��O�������L�B{���\��Ç�ԓ���~��7��SS����*���CK�w�]1�X�s��͕��L���Cױ�.\��LP���Þ���Ui���R�����M��ğS�ֵN�g�oکK��̘��ж��AڊW�{\����K��B���b��


�^U��?��wWޑN,�.�[`>.EY�Ӌ�$���'��C�S6M ���ͧ���#�@_�D���wS�$'m
[�F?q@W�39�Zr�뛝��o_��U��WL��V��^-O3���,-��ګﶗY^>Ї��;���,�u��%ꍤp�����z��yz�'�8�h����â��_k��ը$!�s�O���S7ט��966��f{�����/�x-�wq'������(nܣ#Z���M�E�5�GВ)QS����ᮙ�����h/y0p�Q�IȺz�t��b'���r_���Z��_X��3���}]�QÿӴF��c�;��ޱ'.�#�tu��P����̰�ML|,�b�c��5����p�{i�x����rH)R w�mz���q(�	�ső��������P������-�:=qZ=�[���T�>5�8�-�)y_�BA����8��`#���7�(<�x�V��4�|V7��؝<Y���M	D����Rt�ZZ���n��4xȠ�	���b�H��_f�E��k��L��.s�3�tl���?.�u���a�z�|H���$ 6m`/������u43_5t=
݋���4���O�r��&���`��s1ȰDጧ���~� ^�h�3�u����mΤ�g��y�4R��K�154-�уc���y�n�p���J��Ŏ� b(�{��l������9�#�}9���L��Zf#����D#R���`����p��r�Zf6~uh��7�/���&E���`��.@hy��}/��K��竂����ٴ��.��74�I��7N8�O<N��[|���>��'�y��W��[L�D��ۭ����l�]$� �9@HbD}�2|
��)S���Nܟ��<o�y��cʰ�X�~��W�l�w���n���+4;�k��܀�=d�V���,kA���-���N܏x@zl�6��B�˫��
�ߊK���������g��i�I=���зG�q��n���K���P�575��D]Y"�A+���,�)R�lj�����Z|�,M�N�|����]�魀���N�$ǌ0�7p#n,9�i�Ue�;t¨�3�ܐ*�Gp��q��HF��Wf�J�H�U׳��#�RmF~��4F3c�?B�iq#�[�p��hϔ�{%4�+<���C���Ӏ�婶� 63m��3���G���I.
o��q
$tu��^�ڳV4)�:9�J�M�z�\�d�f�I�˿�be�oi)2=Z�LqM�Z>$�d_/x�'��s#���	�� WKe�������p��feQB�� |��͛ae���&$@���q�>|��U�@~��h���pY��ѿx�A�č�n�]�4��Z��g2튶/3�'��m��y�����ڞ�H@�:W��H�8�-;X�͓jXc=�d�&	
�ΖO��[���Q��y�o�hm����Q �$̾P}g�Z�Gf21����'��G����J�4T@� �2@�_8���n'5��:��g8@9�T�-}]Q6�a�ú���9��!`���"�W%!����4%��8PrßR�r�p�(�&�T���')�+ޙ�u���Ra��7���D/1vm~��C�pF?�h�Ko�V"m����FI�QBC{_��f�B@p+�(��縗f� {��T^�[�7�R]�Ӻ�|!9P�:t���l<썥��"��'���@$K%��E�6�Ѵ_�L,��Z��b8ߏJ͏,�H��bx����������z��O�u��!��MoFC�A�<�*��-���-Q���!�!؄�^�$88����e�F�^������3;��2��"�j�#�h��n! -�6�����Ҙ<�T�&���U�_R��F�Q���I�n�7��Y: ������O�7@z���IP9�B���)�d���v�g��#�ݢ�2����3��g��a�?$KQ���+E&��Hv-��H6���2v�Z\a�����ˍ��ɝU�c}Y����G��%��BuW7��a�����#�B�ӟw���F	�x����i��x�46�Ok�:1[b�\|?���_�)e�2vy�C���v�_��.��~B&��J:�^���o�k�0H�3��Df1\���O���&֢r���s�v5����M�D(E�?���:��o�+B�`G��e��Uw+��R �����v��'�{�Lq�*�qm;ZS2�z�v�G��ޱ|I��i�k��h�/��"_�3�/��.�Ś0�W���h�T���r|��Q���;���D�����{6Jw�-4���S����¡��a�@g�SIؙMx�	����4� �^��Ӧ?EFl���4����V����s8_�SƑ:���7	!hty��]� �z$s2�>{��i��iK݇����'
=����~` Ȁ��;VIL F���V�-��ȿ���P������ˇ��W*s���X���A�>��p�R&׼��,��x���On�d��XPl���͵=꠺�;tKշ�fꞀgh̠Vh-�WЉ'���A�R!*��$���" q#�Ku9��Sb�2�Kc�0�h'�D�j��MG���h�0�
�pI��M@֝k�z��0�3Ҙ��<O��x:�����F�}bk�2;�%����a[��B�=���]`��r}�H�9�׭:s��Au�
�+j��wY��$�-�ftZWȳ�l�l�z"���A\�{m
}��C�&|w�Pv�V+t{\� �v�{x'</��I�bh�'��ۮ�q�����ա�D��w�m��J�8���L� ��ee�R���h�ݽ�Q;�M�0哺T4|�N���c��+�U4�b�,"�ZYJg�n���V��H��Nz�,��$�cx�W��zl���u��*4�c�����v^��� d.9�D���QqOχH�N��N��+rQ���n�����C�����\p�(��G� a������۞�3+h�$�ޱD�?�9���.#�5�����۞fKV,�����o[�U;wI��.���03�4���EE}pYѦ��ވ�Ҡ=������y{�6F9����D��3`��ZK��s���Nh!���k�Mȯ\�#ψ~��̊�:<�* ��e�_�_�@2Q��*%��lΑoS,�4��(55��_�e���P�=R�ϓ�0V�/�A�G�0aM�V]�}���vv�_Ǆ��X]�!�a;|�P�v+f ��*Se#��0��W(�ԟoTi&{<J�����%��2�m����_,Z�{�)��Q]��H�qA����#�4���C�<����`����3�P9��Sf��-2l��U1t��2Oխ��ئ����>�	\���i�1l,�-�G2� z:���K�b�(�g/�ͽ]e�k�V�o����߇�X�5[D*Ĕ�r3l^���ajሗ.2�}��k������*����}�a��]����DG�>A~�i �=��G�l;�s��,݌�\��	��{�d���{�6a��߁g��f�����:���@��6S\2�"c�QU��\�K�Cz����� Z�q\/��}P�R�{#�{�N�}b��\�;pxMN%�Z]U�;�MՔ=Mǵ�T�~�W*���4R�h�@��4Tp��eWC|�Z����̧.	Ե>I
�ys��9(�\��>$S���[t��l�}N�t�lD��1�p�⾖{�i'#b��D!��w��u�ڑ�ܢz����J�Of]i���'�5��.�7��t�1)$$�/���9\b,�Ю�<��R�ͷ�x���32�Ӥ�ě̈s�����3��/P!���Pڽ,,`j�Y����E�Y����ס��r}���3{�C�mz{� �����FQq�&�Bv�Lޚ^�v&jz�;bί��f��s�9�j|���9��j��-�k8��+ڟ'F3����Z�;��O��@�Y�l�8I:�4�`�-}h����(���s����M5�֓�;��UJ�Y�h��_��=�Ϋ��&��z�rɐ�ce�u�I�YO�3��o�p�����&}�&L%ת�ҥm��cL�,nF�� ��rJ�шG�e?}r��@����NL�P�V��}ݓ��U�%z�?�09�e`�]� ���ȿ���t����('k�c=��K�����9^j���O�'�L��v>�}\ڌn����h�y��ٿ$|�gCo�WW���3&�J<}w���߄]1���U>�����TTCe���Qf��C_��^�5�в��L���e��XD���#��c+����$��З���=�����m>d��~"���\lzQ���`����SC��ܕ0��-)��G^ooW�SN�}|�����Aq$�.4��o�'�������T��vy]�p4[n�����.�us��D�E_�C�G�<X���iV��<��C�U.!�@ٰ�7sj�w���)wؽ92�mPr��v��#�p>.Ƞ�snæ<h<�_}�kʂ$W˿��2�!h~����IR>�}�2�$���drа����6xs��Kx�믁�;˟a����2=���%���.N(Z7�7K^��I��RV��A��8XF�����;�:�$9*�宷�x�iqtG����뮛�)��*)��{u�e�9!���!���45�ﾎo��H���bN$n����4�Y���q0�v���A�Z��ס��&J֤�[.��x���V�ߠ�gȮ=ݭ���m@���{H��,+8VX뒞������2I\=dZ�C�.-��giY�<x�W�T{���9�3�*Z��܎om�ѧh]��:�"��;��l�ə��\^��؏}{O!�p����*�y��VQđ�L�����s��t�m�̎s��1q�>GM�+y����F����_847�آN�HR�%���F����D%B�Kd;��2�����`خ���fbe�JY@�q�toL�|��	��j�����p�J�G����o�#d�u���Q���^3Z�@��Ϝ��U\��ncgș�!=p'�@��˂�=1�D� �qK�\���)�@g+͞���;�I�*p���X	?��#Q���f�m2(r��4�|�'�DT�y/����AIթ,��xX�f�`�0��� As�jd0p�H[�cPިe@����Ĥ.���5Ѐ�y
�X`�n�w��*��w8Q��v�^�F�M@���]��R��
���;;]i�E1]��K�n�ȇ���sX�^>oS��5+�]��ӝ�s�
�w4�x�6G��l6楦`�|�[	��V��s3��C�Wj��A��^�=ً���[P@6��Z�1si���ېk_��Am�����65M��6��	�J}ͺĊ���>_|�sL���o{�5��a��,N+�+�^�t��.dj��-���%�C���d�9����Q�F��?�,��/��-�+ۻ�{G{i�"F�J� =��"��і�<����0|A���r���7m��;\>5��l9
]z��&g��7?I��$����JK�s�����.�����it=��F��޽w��{�M.��� �̏;��$ͼ҂O0W�����pE-��2"m�����l \�ں��JW�3�l���هga�8�aE.~������XQ�#�V�Y�v��.,�6^�֕d��)�b�<u>H�,}۝�xf�TY��+��T{7�.��2Y�mw��oy� u>��tjyѫ������tM��#��&���wK0u5�d�D��<_��T2��l�}b���6��]�b���3wl�?��&���m����Q�Ha<��5zHrrv28亡�:|)�
$��:)2ć��t�ŅY	U��G$`�R��c��k�?S黆�RlW��g=��W��fӓ��dҾJ3�Ȝ��͇����L�ȓ��T󋈣��YR���Ǭ�K��F�C%dOS��a�e>QH�8.�|*�uN;*~hD��K��y�+����t�v�^��U{�l}{l���f%�MŅ�*{���c���U�ߊLn�Nz��)���y��#�1����:Ol�nI�Lm��3�G�"
,�i����=\�S�x{u��cJ�b('�q�Y��ug���V&6��1��y�!~�t�o��2����'��z4ݘa�+����\���	��J�vu�1��Nyɨ�xl�If�\�ע��KS�
D"�j;��c��}o�"��C˙�����/{�x���~f�'Mu����L�N�$X��iU"�k6q�in�����d��B�dt������PZp8qߐ�`�+�1R��L��RD��qj����&<����}������nh`eկ!��u�z�
daeW��	-�������(>{":*�ֺ�ʦx������,^	6���~ɴ�'}��	�����I�r�;��p%d#V����/<k�8�W�]Ȑɇ���Ϧe�Ad0%�f�Y ��D������c�*���w:�J�ߤ�*k��{Y-]X0H[�k������x��{�J-
��m�O5^,�:b�M�N�W�����Xi�Y��\����w�K�1� ���ɘ�~RǞ�г�C�\S#��uhE��7�d��F�γ-�b�zHD��[��&,��	�&k9|���N�:��n�cռ?�[�;�  �G��u G՚F>�V'�53�,^`9uR�-�\k@G]�3��Vvamhv�j�w?w�c�av!]B����0��ǚp��O0m������=�4���6���}�|����.�+�tl���z_<uР"�JL�/%���O�]������������xJʱ�����/�A!`�I~�c��0�� )��?��g:��AUV�)b���](���JtK��|xF�iu���|��i�+K�{�K��z�v>|9&(�y�Mw��F3�r椷S�6�fӃ^
=���]��AH�=�]�w��^������ٙ�#?�;��R�ΛWs�-��Z��X��.�e��4	Z���KX5ׁ\f�0�P�'��o�wp.�+��)��p�H�OqZ�ܞ^��o��S����7���})[)�� 띦�՜��u�:��.W�5�㢾���C���Xn?s	J�������d�fއN�Oz�́ۉƈ�6:α�V���c��t�8A|�&:;��^(�䛩8{-˱�X�x|i}�qs.���`~�t	/P�C�ޠ�*kll�&�K���IrY��_��V�*����,�gC*?;|;��$��\[9��g����%w�-3rf��RS�����\����nwWh `�����<jqјzg�;���Z<��3�Bu0�C�=9�.F�#�4����p���۸
�Szj�O���giD���AJ��z���q.;������
��:Vg��T,1�S���e<3c�97W����5�y_w��S¨F�G��c��bC�۱y|un�O�3�/gؘ!���8�A:E����崴�-9�p��-�C��"��;�ɧ�+r�b�O���&ú�E	,�o�	u �z�S�E �'~�n���u0g'���e��Dا�Q��w��a�)7��� rX~&�Ь�?�;�����4�x6���>�It��^�h8�z�RK�y��]�r �vF9�.�%}F1�IL�L���ћ|�_(��\E+v%� V�/���EF{�^AЮ�+wcm�|�~���5����3�V�sl���q�pcJ�).�b��Z�sK$�D�9=� ����U܊�N!K�D��?�������^B/ul+k�o�t�>����c�Y��͒fӗ����������k>�����˱��6�rR�ih�T<���+���T�o�Y;?�tF0XC:��xPC��R���gjs2��e�6�ɒۺ^o|��<��ڻ6ј��L:6����!��X�x~���5L�Ce��V*�m�'����1�nl��;�T"�����LZ�V�H��GQ��<�Ψ�����!��@#4&�r���y	������{'b'�f4rJkн@!�l�Iv  �+v�u�c������2.Jo���iD��k�9Bf�"�CR?rCՁ���n	;�E�Oy�үcz���w���!��z�։!��7�A3F�������y��K��x��l��;�ʐ���"��;��;��r�����~��Ր��f���d|���K[&�Уry�!����^���H�t��2K=I�=���G2wD�e��gg�e�;�G�-]���q��?1��X�����=��%��,9b^Y���9XE2kS?���#��������xI!����	�z��e=��TN�O�*��i@��)��U��c�a�����.&X��%6���æH�[7��V�dn.��U �8	�f	|=���Ϲ��ƪ��gGK���o5�ͫ�}����l�=�U�G�})���f3��k����p����OϾ��L)ra����묁�� ���� b*Ӿ��e�[M>�3�!�aGҤ�JH�#��چ��}�V�ڠ6���#M4��\xAXi�y�����V�*ȭ򘡬���� ʚz��XD��y����S��Vs�4�j��� h�~� w��Ք+c��b��2�����+�_eW,�ښ�g���B<k�^a��?;���3D�k*S���}.G>M��$D�����p�F$`~?;3 `��Y@�7\�[U��^���h�+<�����?��jR(ͦ�x�����	U�Ϙ�\���KM-$�^�o�Z	s	=7�bj/�;��>�k�͕�G�l*�U�r�#0�8�q1T8W���﫩3�xݞq�6��o~`��R%�t�3ᖄ�q�Q8�:����		�,�Z�L�&�����5��?�O��Á���=���WR,�p���be��tX���j g��K�\�U,�#,�f��s��Ba�%���vM�n��ڔTL�I��l*����!9�����P��и}-��8�~��
#��̺�#������sT��ʕM��%��8��NI7�D�����5"��v�coӘ4Xp��7Ph���5/�� �ć���2D(wW�2v[�KX��'�R�x|nm����7JF��)����s����|�y����>F�v��)���uc�klx���z!�Dl7��%-�Uͬe����v��yl��_��b�!TJ|T��.�E��M!b�S���rWO��+7�[�X�~&u�-n���q��6=�4h�<����Z�J��#2�'�	/m���B���oI�Ղ��G�b�����P�I6-�<L�}�*�)�f�@��ɝq`��ƀ��pb��i�աnV�7�f�,�$[��^��j�~@���^�0�#UYqB%X]M�����<ƨt!9�_q���'qrY$�����h���6��<Z�Z~!��e�!�� U���� ��Z��q_�5�{�Z�Hp�3�Y򀩒E�٨o�VGP���8P���[�J[>Mό�hy>i!tcsq��e û�o�iI���IG�n��R����C�U�p��&�*��襤�5^1v*���~vVy@$���/�4
9cT�uP��E��`�Zn%wQZ�B�X�N���ݘn�yX�|�������!�G�~�Ϥ�J�v����ٖ���ia�����E�%<�s�����~��3O�ҙ�v�V;����@�c���+�*�;M�nQV�	W ��5</�C�{�+��sI��V�s������C�S��j�>����T�w�v��f�L[OM���l�lt�*7˧��|���B=�p��}K�{�@�\Q��3��K^vr��|�p�[B".�����*��iU�شp,����%}�&g�N�9�U$����ݿ��z�+*(ڽ?L	G�<� 8��k�6��Su��I'���v��nO��{��YTԚ~D8��~�v�J��˾�������<��[S��iP �r�Q(����I�n!�:1C����V3�`ھ���R���F$����BMണ-����ĩ�;7#�χ�W]�JfM;���يf9��K��/a5�@��6��0	dLE�)M�O���囘Ҡ;�%���d�L�}ir5@�*ܦ^|�78wV���>�>�T����}���g=8Y?���B� �h����v>؆��9���
t���������V�3a![��1f������X�6..�A��J?��D�D�fP�Lw�价������{�u��%���dX�	�[�����Ý)�د-��e�{�ꄄ��b3I(�c7����+��n������a��-O��V���З���+���a���"	�L�@Oo��m!�]�o�^��n�V������E�rZ�UN�F��#N������ύ���CRa���)#]�����˙���=b�����۱��T��Mk���{萺:6�"B=�\��z��@�-1)I��%��|�����z��k��ge��q��qҵ�Gb�{KwW�y���6�qxz�I�I_���k:�tv��N�8U ��N�QլJ>y�z������e���pm|3�ZM��0�S���G�%8�����~a��G�Kv��):TS4<�	p�v�t�1�,�_�-���||�Oq�h{�ϛ�oԯm/�1K5�C6��)��!�Xh@�nT�?�=��_>��i�br��V �_��Yu�A�F�lOSs~��J]�|�ⓁdIm���"[ev�ߞm9�<��gO�S2U��5���KG�7 +	1%�R(���B]��~�-��S�<��G����t
�+$
��b�c\����ռR���AK�̈́n*�󮱵K�H|�Q�Y�s졹�.?�n� �R9��*�Oe9�N_��oB��?����B�Gf��x�'��w�~e$.��Ưlb��7��	^B��
J!�g��.L\xA�2ojatA��%��ʌ�\����i�I��������a`L�yNVtȘj�h��74Lc�O\ nA h�K��x�J��Ç� �D9��V�l'���Q�:�z{�U&�?3:q��W�?,0fA���M�����2�WQ@ֵmtgL6�`Cᮔ�(��� N�H��:�e�4T4�>n����>��F����[�P�A"��N���|�'���2�����wH���ϟ;1����Ӯ�ۛ���Y�g3y������I�� � Q=�[�gHstk��\93V�^s��T$���n�ɘ����
����%($T�#�(FW��F��r����T�-a8]Rs�ӻR:l{kވT�U�l�I�8k�M~ʞ* �~�dn�]��m�O�w�h����gtV��
l�ig]ñ&|��IK,���dM� ��}F����@�UP*ؔ������Sjj���rN���N�d�T��pW�O����*�5��c�â����QDP@JAR	�F��Α����D���ib�!��$��;��<�������>g����^{o�K�/ ��p�n�&#��;�V]w�����n�T�n��S��7�M�J�H5������նGo.1Z���?�C����~9_�:�TM-�d�H��$�m}�[J��
�z�Id�L��h��ni\s��d露 �m�.&��8Q�>��7����h�ꃜmY���C�����ӏ{xU��)Ȳ�I{E�󉽺��L�� QL�XwWn���F-�\�o�4K����2c��Z�5�i�,�T�kڳXJ1��F�C�[�&��C����֛��+�
�	��y}%�<t����k�R\\�^&b�0�v9�p��^� _��̒��KXf�[��a�.w�5k܎%O+y//�l�;�m�޵�"�U���W�FtJ)\��3��I��R �,	f���i��mޏ5��z)���t�Ҿ�����"&l�z�:5�\�(*�`�W�F����T?�SQx��Ӿyg@T��t�<.�l�dw�6I�+��:J'�۫�S�V�#����t����Ώ\�݁�o���&m�h����ó큣o��ioI^8"ޠ�q���#erfhRV�[K7u�v�H	�&��7a��j���lMJ~������y��̾�o=%A��q�]�^%�*�> �65=wy����SX|�f��=M/Î�-՜�@Hǟ�S�����ѣh���+�~&�g��~a����L�l'�����Z�L;�I�M54w���f���W�u<�Ϧ�t���pG�DW��o\x?�B�bO|��^J$����t}��4D���d�~�[�D�O����M�+��ۺr U��T���B-3���؎퇣g����۸�j����,`~��*�a�C�W����}���M�C �e��E��Tu��q~���W��v�A�I/̫P4���x���u�[o��K'��d�mC�����[X�NKb��V�_]�r��F��Q���1��cY�����Z4��8�/'��8�0����-Ѫ=DgMX��s������Pw��)@��"�Ï�؆�O��Ɔ*U958'[��o1�7*s�rbп�/��ر����Ľ#⟬8ԍ"ӝ:�_�����h$�u���ER������Z��^:'��}Ӟ��~�������[�7MI������y��n�����e��;r��F[����D+9ܓZ�FW+�b���^V�ֱ���|�8���>�z�k.�:΢�b��2�0i�;���H.�'�
-'v�N�j��Ή!�W��dw�����1�w|��-�����D%r�o���dp��_�'9�'�����"�M',8~iZ�,N�FQ-��w ��h�� �0X+�
ƥc���)�^$��N��l2���߸�������Jg�H-�9��#��i���~_�F����f������e	Q��v�ʭ�mh�r�5�3���EC���{�a�gktk��=�-�����L݂�`	�[5m���t�'e1�����l�F�*b������dJ���a�=-��M�Z}��2r輰��|�nw�Y�py���&>}��x�m��%����Al�B��z�O���t�L�B����i�nOm�Ƴx)��o@<BZ�3l�g�K�����W�򎄋O���G���� Q��5�਱C^����X?@���΅&�	�j�-"��C�m���t�FI�
�ĪK�͵�$ej������F����)��<U&��^�%SL�$��\�=���^֠�D�-�]�Xţ"-m���3��S�bه���G�8Ḽ�S�r����lި?;:b��7�.ǔz���3ti۔��?��=P7�}&n"�{fjPk�ݢ�\�E�v-i{�r�G�I��	���W��-�c�Ddp���^{�R�&]u���ˎ�K�!#<��Hɑ�-Ȓ�Ї�WuI�5��~z�f)ξ���� ȵ��n��I�/�/�K%'�ҕ%R�O-���a�+o���ŋ�h�ܱ��o~!���R�r(����h�y�S�{��b�P��+	f��Dv o��c��OW�qv�Ep\��[g�j���+�EF>���}��*��n�5�ۧwg���rw�>C:�VG�w']�F�ւ8Լ���� ��y張%���cn�2��F���@NA[�w"N5f҄_ԶT��,Mz{G2�-[���9�m^_l7z�{��.Q����g�+��̭��y�nL��Vх3��֧�9@���d0Mi�w��3��$گ�LH�d+Kˁ4L�g_J�}�4�˭pM�
����e緧�dBX\hr���u��"� ��Px�[j����6�R�7K@�2z��ܐ�l���Aa߳WEפyM��||����s��y��,�`.���H`�a;���&?R͸tOa�!,���6,�6�8�L�{�;�K�����o����U��c��$SY��}O���˩`�AR�{�������q15��W�H�J�Y�)j8Ơif	�ʅ�	�b>x�Y�P}T��֠CrG�Ϛu��~����qLx�,���
��}����v�j`�`Ũ[��G��qQ�ب`z��uӄ8����{e�@�K��]�.���M�����mvw�T8��SDJ=�I���xϷ�o�;����}�.4�|d�R�|�#L�:ܞ�(r�[�� �V$���g[���� �d�̽�W��d7@���4N~�|��&Цg6�A2PC6��� �q=#���E��� ����8��7��,Iz�>����q��X�t����/�T�1����I��Zf1�s�/�~����d�:���4���a�h�Sy�����Iyw�Mx}�U)Mf��Y�ԥ�?쭣�N�˕N#��v�/<Zo
����LoDtQ�p���X�QC|���ŷ�H�rJM~��#�;ـ}H�fJ��M�6����:&7þ���&���!(�n���������U��CR����h�O(-�r`���o��c�V�����D�өF��%�D�ʈl���n�s
cA	��6��8��:8�F�ܯ0�߱�q��!!�'-�wah�c��J��j��VV5�D᳐s���K��#A���=E��7��̻�7���-�$-��<;��w">�t�s'�	�q9����|��ӭ!�-���\c�']U��eG�pPs��\72�����N�P��I�v�����m$��k�|�_��G�T���TD*��*ؽ�0��T�JY_Zx�����:���j�L7��(�scaQ��k9Osvq!'����;<����.�m��fa
K�����)���C1B-���	ub|�p)X�hC��9Ŀ�r�8��`�j/g�����ظ\���s�Ol4������E����
��=��2��E8�Y:�cU8�&(�LK<�9���n7n�uç��X6�� �/�z����I=�`D�?/�]R�AOH+�օ!JyCe~�@���U�/0�Jd8p�Kg<<���Ϗݷ��ĽV"�>��J����&�L��Aiâ�gK���Oy{-I�	�w**��%i8��r_��Ⱦ8���K������tk)JGz�%:��۬C^�2��(h�U��kLh,��eY���ي0� �~��8\�dW�/Z��%���^s���~=,��(G����VUJ#{.�n�#;HZ���,�mt�	Δ�}q�I����3�@@�������}���Z�E wk^���2�H{��]W�6��iy�O�9��p���oZ)��-��ǵfP?�<n�տ]�$s#�Ȯ��q0�(�u�'�|����щz	x�j�)��x�x��S�?vj ������{d�Q��Sd�c6��x@_��Mg�	E�TZ%�~EeO��/d ���s�l@6fLa��������P̹G`�5����+l�B��0�/�B�߫1�VC\�ȸJe5|���)��faҲ�9a�S��\�*��F�JUW�e����9N�����$x�ӌ���%U��c��
��0�Y�����y&#���X�=['Bt��H'�-jf��4zI���f[�W[)���������U~�Y5�Fn�����#w)��C�B�Q���A3�h�|?8�%������ݽaӐ�K�?t�&Z��G�&�4W<����g�}a���@u� B�]EcjLC�C����H�D�R�+n��{�\���:E��9�m嬥&��!�Z��<�[u�{����$��}�Z�
�P��a�K�%��Z^�*��\V��/,`������z{ �����=����n�j����=�)�%�M��Vur�z1Kәrq��Y�OxĵR�!|7�'�� ց7�".~��T���-�$�;{�ȣ:d�`5z��h��MP��_�g��"$�U�X�S/�n�=^��j��j%�/��o�c�v�뼸4Nƒ)+=�E�A=��ba��|H��BM�Z�e�53d��S>�\ż���S�^�9Sw���#7��=%�F�<Q<aoۗ0�[2d@�M�$$4v"ė���k��R P�tϟ��ꁸ$_Z7��i���^h�k�nX�����I�I]������Ȼ��ֈ�ɰ_�;Y6��n�ʻ3����	\n����������1�\�e�Jq~���jB+�D���"{��
W���J��s��/������W�qBGme�Q��7W���u�Dp������p�Zf�P�N@y��3GY��A.q��T��q�%�����BM�]��j��ϫ�,�Y�F9�~v�y��l:4�M�t�b��_�=�(%������}`�������(�����T��q��2����G/��1��Wn��L'���jz�_�b�(9��3���/hH��q+�;Qx$J��O�&,\���Q��Ҩa��>����v��̢ח�s�:D��}D�x����.B%����l�Q}C{ ��d��C9����7A���K��8�)�z|
��)��d6�ۈ4�s��r���Y��ဓ�23����
9�3� b/��ǅ�1���l(��A�7�����L�F����k��z;��/Gg�x̣��?cbW��r���,zEkz��I��px/��]�5�$zM�F%� ����s�A���2���ez}ݜX{m��K(\���?�0�'�}�f.29��.\8��U�\=c4ut�T�c�0j��x����X��U��
��=�AT�@���c���[��"ݬ��M�0T�4b���]I^�K�nS�?�0���cN���a4V\ӏkT��UŖ�oЂ��㷍����,�����S��=ψ�r�N/#9'����3Z����d5�I��
���W���[?��PXC{�:r,a�R����"�Na3yQum�{�b�\�)�B�x9�z,=7�T7�KNp�JDbb��b�x�洰�����vD�#���B�V�8�6�À��[a� I�kq����;k�gQ���ۏىhO���;��:��ɨĿ�S+��`àQ@*�ߚ�EtǗF���n����{L�AD���[a��"�o	O[�/ �o�9����	��A�f����d���+?#_t��fqn������g�Ʊ٬%9O$��*�u���[-L�*]� �d�H��"!b��3�C��먿zZ�ڮ �3�V׼Jţ11/?.jjD���B�z����=
�4+*rn(4Ϸ�d6�7�����K`+u���������F��&pw-3�;R�f��i�H���瘠[hb�@�q��G�&�:�_:�� 
�{��(XQ7=L��<&�m3È=UԙQ�DY(#��CZ?�ƛ��Q�I���]w��A��g]A&���_y���;"P���)�N:6쟫�$g�S�,*'��f"Ӎ���l���sԩy��̪)n�{k3�2�-���x6��B����Jn:
��k�55/�R��0@8���ۨH��/KT����>d��ցd� \�@?��n�o��V�'
x�Tg�5J�M�<N�QAw�\\�De���=�N'VM~�A梪C����a�c�@x.�##�w�9U@/}���j6�q������Q���o:�n����ϕ3Jh(TѰإ��U�C�W��n7�/�Iٽ��M-3B�(�?��O�R~,O+Q g�����ǺĪ�j.BH�/x��x	�(����k �����ez�Ż�q�Vl.���K������-f���̰�k�:�Đ���� @#q�/`(�РRL;q�ϳӚ���
�_\2�����ql�B�:	�:�d���y�G�U����H�C4����ʸ3�4��ޗ��7f���<�T���r�Qj0@�����6((����Z����h�3J�i�Uv�6c3;O�Q��ɒq�h�<!�ʿ�:�G�i��M�����u�W6:d�Y�D�:���"�)���TCkh Uf��)�"XpE0z�q,�lѓ�J� ��`�Jퟨۿ���L
 �1��w��eg���#nf���J~�H���5*G����i6"d�}B������
3U���K����6��,'7Ξ�F�������rO�����?!Ψ�N&���k�-�U6�<��h�O_W,�0~EŽeE^_{��C*i��A�`�Iw������z1G�>$wjQ
6����g���@�}p)y�{�5������k�A���{@���?����d��`��۾jf���{�A�V� `<��2^�r�Jλְcf {�v⿿?y�Qs�'x�}5�Zd��sv>�=+��uG����Z��p����� ���ì�	�s�{'I	�le$���/Dgss�"2*WO32�/���y�l*�lIX��a_o|<���I-SG�K9_���Te�l�](C�a�l���v�lآ,s	�~U�=_%� = � ���uӾ���Ռ��f�$Ѵ��#C-^��"�p0�*��X�Y<�LK6���v|r���ĸE���y�}���%�t� �a��l������0`P�d(���O��q�)o��t"�<�q:����A2 @Otl����ChG%�&���=����:���VI��}����|4���৭Swf���R�(�-�T&O%.�z��쏩�
B���� �~i��0�>����	� h����N�N��Q�&8+H*j �!Q� �^�� Ӝz�j ���\�5�rQ��'!��7A�'.C�{L=�.\������ ��K�Jw�aR*��ڍ�-�<�!S~깚<D���a��O�� �p�-�a]���g�L+�G�wq9�%���߲!z���ZX��sjX0x�A��B`$0Z���`&�R�p��e������c/̆K#���gL�m�ŇUh��\���s�ل�S/���x
h�R|�T9�9�~ݔ1k�p��D��OU�����m�A��m��e���G���w������0+�z�ߠ����O��Fr�����5w�t����\��W�D����[��@|���JU��:<{�O5��墎~Ң��~z�o-|"�@��D�z�{�@��X���u3���&1 �@���L�H]�ss������	Q�v9{Vx�f���;4qh��Xb�� 8ė��G�'QA�4Y���B\�B˱H�},*�\�?�b�v�� �ӻ���c��w�6��4���H�s7����_���s����� �x�0�Q?5t�#;����X�,p��q9/w ��$�Yp���:���7�M>?᧏�������&�mq��h���K�Lm�/;?O���-;��,��c֯R��[W�)�� �+��4 �䀦D�B�9;b���)�w���oQ�ZP_��� b-9���p:����r�Q��\z3�N����r��t9n�q�����q�@/-��J8��9��U�^G���5}tGt��i� �ϳ��&��������;k^ir�$;G�ql�^������Ա��϶��(�h�f�!'6H��� �0�o�%��/G2���r��쥓@|�8:�KVSS�Xdt8;6�.���f�M���f����#��^��{�a�������.��X�?�cz���CyrpT��>�{�K9: ���kArQz�����"2A,�|�;W@���7�`&�)�>^����9.H��d���v\l[]^V��i��@� &
-yӿS�-hי����R�'3B@?���m���kU��0&�X���h�BN�1O; ��B��"2�2/�l���z����H�O�z��0a�i2�7_3d��Ц�B�w�2�2��Zeӄ������C	E�
��^����~s�'�l"�t����F�m����$ZQ�����"�r�F�k.=��<y���Ta�|g�^�ċ��銶��q�W8�=�P ���Dk7�Ϝf��z��V���)���i�]7�O�s[�]�r X|@����D�o�	`ܤ��8�ߥ ���������n����sv@ԧ'��j	����皵��d�����{�:M��|/%�6�O�M�b������7�m���܉�%_ڟ�6��-A<u�^�v-f���Н)̲[��~�P�������#���Ωaӄn(�ڽ��%cO(��b�����w�s\�0��9)�i����[�=������	��!읃:#Rn��ƽT���$�h��K���VbJnx��4�n�9��[]x��I 翽08ts�}e��O{)�%L�#W���o�R�o�D᫏O��HG��;/�8>�J�e�1��[�h
fҤ�:��Q�6m�����y��J���N���}��2r�#�ź;)B�/�£�����U,��͏Ҭ���A�����}��Rx��P;���٬i_���.7>���qM�z�0�ۣ��6�؝�x��(�|'n�\p��+�
��| ��S�Jm����Em֎�dg�g�E*���i�v��S�tM������������TQ%`ذ^/�--�^-�0j�qSD��Ɛ��]���F�/���K{yy�p#Xg�'s�U!S�`���	����qs�W���|�c9gꕡ<pf��ڱ�<{-��|�s1�9V<u/��{��݃K�TE��e:1Ҭ3�����É�����ł�o6D�����Π�����rb�͇�-����#`�>Y*�:�����v���{����Qk:81.�G�)dI��&�������U=��!H����J*�,Ü�Z�d��U�]tGn�`�qu�K�~:^3(�iK��hy%�?Z�%�����t��8Ё��/�(���Q�*6�,�u��1�m}-r�C1��y�|�X�\��k��HK���ޭe�{��.E��B��䗛�J�5���I�`M��
�z���j��YCi������>#��
1�u�H�@k�TWjfc!d ^���2�6���]���",��#0/4��KR�	~���fӽ���dcj��%�J>$����(oz�R���$}�U ;_�r�ޛ*t#^�<�ՂLik��3���S&�E�%�:��X̼��w>ꜰ��>A��B�恛t�3�~ᠹ�I�g�`,N�	+1�B��;�i�T�C��6/9*M�`�b�OL��� �z/o�?!�)�:�q�EY��Ch���\���4���F�@*9<�x9��@�����n���ݞ��ڳ�Q�"��.�j}�- �&�>�����cPg��s2��nH���M3�~l<�������\�::�"#�*��IH��������q�WᲑl���~���"��e��ly��+�$��g�nOҖܐ��~=�q�	Mѭ¾*۳�%�\lӭ>(��-��ĸf^]*���wŦA�u�lb�1�$�U�M�"ϻB
�LHDӷ����KQ��:�8�~��R�/E���m���r��.3<�Z�w�o��~7�(��v�C�5L�=	�^i�G�HdK��,s���������w���A�"��O_`���՜ ��n��j׸���&o�>��0�%t���vUS�s1���ɆM��Ns�[Oas�Jd�8�������l;'v
e�������6�<x����α��rO|�Ǿ�}	��W/oMߪ�qB�
���)l�SE8S0@�*k�����!4��ߚ��/�
bk�>���/	�����
S~Bq+QΏ�kE,�~���x�b�f�M|!���e並}�g����uS�Fop�N��T{oT����-`A��(�"lvFnT�0�؟�w�}}K��
���h�]�̽�׎1W/;<E��Vⵖ�t۹E؄�����)�E�&f�Pg�����[��zN�~1�q�b.��"j������?SX%f7����.���N��m�W({�^ܕYgCkP/B(?�J#�3<uB���&��E�ر���̔��,�nՙ�z~��K~F[����;�Ćy@���������� �K�hBn��s��=e�{FB$���l�x������B�,�%0( d�z�I�������(��n�(�,�ƹ���[Se�V�^l�k'^|[oӵuR��8��6�1u��]���(�(�o���c5H�=E���i�k;�G�����hX(��7c�X@_���Y�($����u�#OA��[�� �����+E�n\�A�Y���{|C�'�����%���O��NLM̨��C�d>���hS��4= �X��E����gr��IU�,8�������ոK���h%	Wo�%����j��Y}5�l�ҶU��>v�7�e�.C�J#9�F���R��j�������!�8v��CW9�kW-�%� �>{�b&q��#%�I[��6�uq�e;tLj��,�����m�·N�~��=^�
4o����X�hJ��Q�6z󚝪�FxĴ�p��
,�٧��t�F{�o�.K��b�T�Z��K��l��*D9�:�K���.AdQ�w������ ��H!M�C�<Ϥ���d(��+��>�^Bn8 z�_M��n�\�t�dp��!���)��qa�8��Q�]�a]4SV{} c�9<���*�X�j�����$�tp)L믅/�����^ h
�Nɟ����C*�u�X�Ĝ���{u�
o��;��5T��[��ҏ��4V�
2j2䪑	��eF^:�~�.�?�s�x0��=��௪�Kq	�H��(;:y��h첋E؈E?E�=����Ƿτ�ƫ�.65�	����\��Ĝ�y6��6�O;M�u-��ع�K)�b��u����g��U~7Fz�[�W"��z��5��|��\���#��2�������Ї�x
��6m)�����z���Z�O���,q��g���FP��iy��%
jګ�.�My��7����b��k�/�ٗ�Z��65g��xe�t��ce޹y7�j7�p�H�^�@�TE�ի���<��@���֠:��r�V�^m7`��*j��%�_%.O ��7QU�+T]�r@�IT�A��SH�MI}7Y������LY)&�!k�,���W2Qa�U�0�ח(R�8���*M=�ч�Wȣ��NZ�<W��#�b���)]� J�����`����z3�WϠ�����]����d���x��G����*jF�6fgU$#Pd_DΛ��%��J�`��L��Dm����~�����z����b����ߜ�R��z�駋Ҥ�K����xصǼ��������ݣ�R�Fj�NWغ�r�uu^��p�=��_ٞ�7;�/�*1_�<�8<��{�0Tѩ��;Z���<�p���K�����q��r	������Ӑ^�YA�<%
���ң�I�K1�����aw�w����۝�+qPz���f�
k��i���Nj���=�)�-����(����B�{rÖ+a�p���%ቻ�&>r����U�l|��r
�y�*U����bN��T�'�bi�%Fi��Dl`����gowA~i���$��QG�͵_��r�Ʉ�2�dj��H�{��VXI�,��N�6�u-'��0����4���SXEe�X��R�m�\]sZq%����R�,?��𕙖;�[�7`R9�������h� w�L�m""}�mu��I.g��FߨhQ��rbP�����}%|a��9���H��q�c�D�U�n��M�>L����Q|���ܥ��D�vMc��#7�9�ر�Jg�ǋ�&��~����)G~�O��<�\����T���0jz���9��eӺ�s5i(H��������m�;��7Y��d���إP�8S�;9e�7O�{>�d2T�SP���{Y��>��~��c�{C3aoN��x?J�Q}�pJ#a0Y��Ļq�h���������+�3�`����T��9�݂z�{s��=��ݕ���ν:����~�S�,�Sg_�6��W��.���o�&ANL��Og�WË��YIoOlPT;ΝN�+�N������6���,���V�Uk$;l�Kc��A`&��B)f"�;��_6�s ��/�>Y01!!fb�^���T��o���r������~�kL���t��Oh2��jM�	�	��Tv��{�|C��};��U��]i�CZ��2-Y�ЊT}̴r'�>P��K�� 7Ks�3�ۻ�z�\*&o�vn���(�H�#!��+��C�ƥ���yX-�!�_�e0#���F�2-�jEg�TR>����\B�S0,3�Y�%�.jr�4�����3�/ߍ��:��Ys��s�}�H7gi������4� �^m�;ݦ�",�ư�xd�s������[�̀Rx�� l��� ��`\�n�aK��Si��N��)�V����V<���o'��v��<�l%M��!e?���)sΎ1��4�o�Dp���"k9եlɿD�bL�� X�,1�~	��/��u�;t���(�H����7��Lw.�������y���18YhTŠyA}�9��7����)�;t�!�K�$3ˉD�;���(*ݚ_q
;��6'd��Z�l�Nˉ2Y���}�i�����Z~����K�
�8Kq;�(��E~v�=���Nx
�/ߝ�����7)xރeV@���) c���S����g���iyt�)�k���PǗ��gd%����GIK+`%d;o%WD@5���N�b���7�7��Z��w\��T���O��P��f�붰��M�d%Ak׃f�Ղ�������n�b
#ʣ������&�����#� ����9V��2��/܆Z������;�#���r��F����%��-��^{Xx�1D����:$����Bl�
Mi��N��i:p��SL��?L9���S]� �40`n8}�I��ס�bz*��Г�t�q��r(r],�_��i�*nn�],������M%̓�����4���T2B5ۋy���0��Pn��xKôzK35/|�k��	58�Y��&Ll���t=�X���ae+��ث�չ�-@v�~� ��D۩S��P�/? $�/}o������p�u��+땹��D��2�h�C��zb����c����m���nn�����3��q�IF�Bc���ʽ��2>��0ެL��WY5 ���(K&��c�`������v�m0:�i�`�7_Z��������e�t��Tqp|Z8U�Ʊ�b��=٤�δC0�TCW�NFK{wL�k���zțVq���F�%�O�s�H�/���?s*�;�a�m��;-b����7�-
�>�J [6Ј�k�#ܶ@��M���T�*����x�2Zwo�y>��S)��k ��59��u߸4�Wة��.`�u�2c���p3B8�w��j������zy���/��2��j�O�I�T�/A�E�e����f)����^ d�
M��	�1	�U�����g���]|�����	Q�����8�"���������V��p��r �ma_�ի�u)
n<�U�i��>����y�ST������-OQ�ǟ�FĀ�����o�ޱ/z���*�|���,��R~=�*]%)���7��`ms;���]�hUخt]Z�p��~
ݪ��L>�S$7J ��m�.��ꧩ�?��_~}��3��Gm�LT�*�����9�m j2��3�]{�ZNɭ������p9oD���x"M�C�*�1��\��N���������Ti�R��p����')+!�O5n���#�h����:��q�!W\�0Fj��M�>(ox8�m1�>C�!|�ޕ��$i���b��k����5�jH��$S�C���\��C° �%�) ��5��S�4�R�\�IF�W3Er_	�{<������Wai�����D�q�X?��s]8g��vr��a˗jT�up���S{		+O��J��Om�6���������/;^�Yg�o�2����&�z����%���(�P[�i�4T�N�t"��5"��P��k#���յu�א��}YW�R�.Ԛk�]��V��3?6lS��ymN$�:��S���S32�)1f��ĖY�Le�|�"����$��
*���n�����Ig�3���[��L���s�(�#��1��R|Dҋ�KM�8�&��hKـ/j�P�n-;���P����@ˉOo��x��;��s���u���D���iK�|�_Z&>�n��!"U�/!Zp�̡^R������n��EGB诳~#�t�ۼ�ڞ���3
��)Ӟ'��f��y�u(�J�s�7�b�W�|uʾMx!��spl��+�ow ����D䖯�$"�@(�]�Ԫ�y�����)+��V����k��G��V��[�>�O�x~�7l�f �x���6d��ַ��Oqͦ� B�M9�A�&�F�U��V@���Smw@��uF�$�[�QE�m����d����S��3M�C@����A$�YW{-c����R�4�S������b��>EB���9g�%�;�"b ��m>^K'��B{9Sތ�r,�����d�0?)��Q�������XIp�B|} ��ޝ��t�D�bC�O.�~B6Hb8��C�&=��F^Nt.���Ꮗ�L�˻�\�=�S��ʫ_�c�����v�J���0 ��u8���s� J���;V���
�+Hx��'�/���u����a[�dr�
q8�#�$�f�C���#MB
~��:;�'�&�����A�i��pջ����C=�=���;�.A������9�z��r$u-W��Ia[2�h���x�-.�V/WYX�H!���A�@x��Q�HE"вQ0pe�~�J��-Qk Yg_�ۣ�'z��')�Dd�E�k��4�X!����o�)�����:���5��mG�H��
{1�]
�d$����{�9��Z���X����D Xm�T{2��y��$�F�䛦�JL�t�q!�r�l��!��y߯�&y,;�I���K{#��S"ױ�S񈭻10��Fw7�\�q�P3ul+k�>g����a��ѓ*j'[rmlw�.`ت�G�1�%l��6�w�#�a�Gh,G�������[)@?+~%�����c"˷�ֈ�,�j��
�7�f��s5ﬖj?�����Y	-���k;��-`0<�K�>b���N6tP�foE�ܡ/�?-���{u@���hI��p��٣j�*�Vm��S[b�4�i�����Qe��A�7��(P'y/g X���Y'D7���R��}�Q!"��I�;�����fZ��$�	9���d���NH2�&V9�˅2���V����m#�
��;��GKߛ��1�7	�}y4��J-1���K�x���?���_=��^�3�ƭ�K�K?z��!��I�F���ѕ�4�o<�:��^��4Xщ��b�W��ӄ_f�v@j��9�G�@�����l�ߺ�	������ߴ5�Ba�e�T���f�D}��ʑ�۞g���/���y��IW�Z�&1�:􍒧2�̟ӄJ_��e�gs����{�!I�x���=��a��l)jj����C��e��o�a]c�܂�����$�����j>I+��r�^�T���'~h>7WןK�Ap�S�AA����2
���+�� `��� ��i}� 'g��6@\��8}�?Z�����W{�aj���<{-`Df^:��ߗ��GI��	�q����OwcQa�%%%�G�?pk���B}����'

t�cQ��ז^म/�I�����	�X�2}��k6`i��e���l3
^Y�u���J�0j�G}��ԣe�|�轞K�Ӓ���T�[���H�kk&A>>A���'����l��m�xd��]6���D/`$]���82�Ȃ��-�_�90Q	L�,#o�1!F�		��4�r4���jjTk �B z��G�<�m�p]]~018�K#{z0�wv��b(��>*� ��3�z���D�K^�LN�u���L��%Ɠ���6���_������w��ō�������Pw�,we�M�dX%����ꞆZw�: U��c����ߍ j�6g�V
�06W8N�Ե��EQ������{�ը�z��6�._B�l����<) ��-��VV��$w��y�<=�xEY��"/wq����?�ћ���S].L�s���E�ҳLt�m�s��]���cO����DH FG�L�/�`*t�+Ͼ6ӑNf9Qa�P��2v1�E�����������un|��,�{˫K�ʦ?�(���C�=w�Oeeè+p����D�Pp�O������%����ܢu���Q\��#�h����qP��H'�I)����F�F�,�[w�:�����s亞�?Q?G���:�˝����9fy�h��n��ν�n0�+ܓ�����ɃN����l�V�_��dؽ��'��G�U�wCTB}��e��6�9ń�I�E�J����;o�c�%l���Tm��y��!u�Ն��e4��ղ���|o�=iȓΕ���QQC��Y����I�o�c�>��a܈wݳ�N�:&|n/��a���#%����P�ۂ"k���x��:/�\��|����������Gs^�)땼��[u�)j�FM�h9Z��(���|�������!i�$�i���B�˙d�Ϩ�X�X�g����_T�9�^ڒO��!�Zt�v��Ǜ6��������ݧ�V/S�Z睔
G\�F��J��9�*ԏ�Z�i�fo�Ϝ:>���F;w�u�<��a��K���c�{���T�6!���e�������\U^�G�+T�
���S	��ieͧټ�aŧ\n���W�u��'�Ss���7��SP����ω|���̩b��������lP�t��-��S��7����gf��|6Hrf��a4�/�)V�9Z�!go�Ÿ�1nf���G��-=�0��p1^��A��к��`<O	w�O������r.�MÖ��0%���=���*��Wݵ���u�̘��Sՙ��Eg�EQTQI#3c��S�VQ���UA!�C�ִ��S�,�:$J	��S�cJ)I	�s��I��y�6ϟ�~���k�����}�}�{���v�W���z���������<Y�-(�-j"~��!����R����4�s׍Ĩ%��aH��t�|�i�7��7塜?��m���a֥��9�Iڎ���]9��������v���;Hj&����Z�.mg��W�_�!�/RXt�L��'�[��k�m��ͤ��S�����"f�ػ��ɲ���o~����3 �K��������x^�W;��->��X��ן���6���ȝ_�rӄ�-I3ȅH���=Ц[p���6§ݦ����r��q���>>g��[���a%��(���j�;��qX�Ґ.�׳ܘ��̳$ڠ�s��J�ݤ⥖&ޮ�[U�'��G�_���"t3��Z[�3GFY�[s�	��#�۵����G�L���^�Ll	�V�骴�ڞ�z�:&��O�n0e�5��y=���t�+z�{X�{#<��~F��l�c&ux-U\��k��N��.�}TgC�h��� G�[5�x���r ���D3bc��4B�.�>�0�b��4H(�?�I��-��臢:H/���$�f���&�1؍F��4|��.xt
6H�����՗�](�.�#����,�y�(N�]�c箾Nd��i��U-zB����&@���*�(K���2Vs��K�z�Fٽ����֝C!w�_��m`8��E��3�ؙ�ם,��#87�)�>+�4*N�~�@�g��-�KMe�r3gֈ3����T����Ń�?[��*ئ8�ʪz[�x���z���DK|�|��ı�;�����w��q3=�R�K٥�ՑRL��I��q;Oڔ�L��6���Z.6@�k��{PjH�Hj'��s��'^�L��s��j�>s�U��Z�/�X����j{�*�6S���@6���/
�L�&2f=͡�u�M�P�E�.a'������'0� @u����s���M>�k����L����H�.���TKnEQ14ec���r"�� ��8gd�y7��ykkw���0lΙ��7��~ct[8�&,�59m4��S[�Ȁc�n��K6�-3>�ٻ�|ҋgEԣ�I���������0 ]Ac�Y�и2�c�\n��@��^ ]׀jn�W�$ϓ���Z�5��e�1����)h%��d��$�������Xo4*��k��N���N4�U�7|�H��tȗ�}���|�p,ь�~���z��;|��]����+8��		8a`�L�EQH5�:
;�`���?+^.���<�R��~���x'�=��~a`>��Y	�i-O���lPE}Vw{eV0;�j48�f��A0�l���l�k���?O?0�؝Ѳx�|�{��\��ނ�<ؙ����?���4�q��a����V�Z
���a���N$�%��Q:��~Vl�����l_8�=<�r+���U�]P�����e�c���|Fvc���v�hb������2g]��s�`�>�S�$����W�{_KcU@��fǄ����9Ƴ�jG�I��l?� �qi�X��C��Wϱ:!���V=]��7|Do�0y�|ͳ|5��HI�X8Ӱ8�=O�G����2�a�����m���������b�Hst��vIb�Ѳ�9�C��'w�'�P1�̘�R��rm�٭�<�
'DK��	>IIYY���Gh`jC	��ղVI\����H����<~Y���4��`�w�]!�t
vس�%��N=�zS�����I���e��k��hci׷�bI
���$��z�XӞ��:5̠k��G�U.UѰ�hW���۬�q3�������n���h�{��33җ�I�W)]��?���5P���)�D3�Y�a�W��@O/3K<�������s�x��j�g����6���NL��E���2�U�\��<�k Wm�q�#�>�(:�ҍ
=Shs���l8+Y3�m�ź�+͖7��NS(`�D19O3������u��Rw&���Ly�� b{َ9/R�C/ۓ��)��e����EV�^f��� y7GP�R�3�!��"��F�1�q-S�K�ǩ�����I���0`����g�e�E��ɝ_��?-FI���ŅzkD;l�f�x��D���j�!����4��`�I��L��fRX�^ї~���[x7}���-D��]�Vr컣�	mL�[Ɓq�5�V\��j�/z��#�⸁6��O�X�RS4Kp����m�|�C�5��/W֏�����fZ��v߼f��OVG�>�"�5�i`��ͷ�`s��8P�)>���VS]�*����|�y�94��Hz��w�ݐ���	M�ݍ�w�>9P�'�22�g_Z��||�	(?4n����1�A=��M��{���b_�����cBӳ�h�N�폯g?�+%��Y��G)�D��xC/�PA�e�C���	���`C<��H[K)(��H�OٜX�S{�S��~1�FW=�IƯR�E�lg JZ�0��% �+i�koL���G�</Q�0zy��5Ѵ_�b�9jf�5ð�L�o�n~�o��c�߰��z"rs]��3,�mZ:7�������Fq�M����#J�gg8k���={-e��0�C�f�Q�[�'�$_��\>H�v{��0������\���!����S��\��*��Z�S�?@:�jm�L�0 U��ȯ�{��P�t�V-�T1ڟ���Zp�l�W�(b�&Wc�����0.g��Z���dӼñ�ѽ���ʮ�F��;�=��r�T��P��Ǚ���
c1x@a��$I�+3AϏq�ځo�z��Oy�\�:��@�ژ���
 0����mG�1���"S7����x�],єA �W��3�f�a�xA�j�0yB��k�^������2�V�x�	]�����
��`�+�� _��E8��&�΄��-\��+������S$�l��d�t#�
F]�^�k��	!�X[�V&�[�PwJ�vCc��D�o5r������]P~��cd��\Ei�}��.�G�
�D�c�~A�gD�����^�X�r��~N�k0�M�KH��o��"1��iIĥ8�P��P��'\���z���Y����/�A?_�*�6jg�l����Z~���>J��0��҄{�����A��r�E
��������;u�kR�b��c�r}�8债"h3��|�դ�r��⢦�z�:����PU�6_t4q�sҫ����!LSt��+��#�Z���� �������_�;U���!T}�ϸ�2�,�R!?�0���M��<w���³T瀋�.���Ҭ�QC�6g����|��h�F�gSs3P��G��e��e���AD��e�х��%XV�tq��̑�n]���o:._�tw�X鍛ԏ��9���I_��-��#�}�Fk4��F2����m���N�p�����F�\��_���3�;�vF<$�8z�*��K�$�����?`l�\�`R�nn�t�zY�4��aN@��B�r㬵�j5ƪ,�Z�_+�a��{�s�N='�c�gE��F�mKH�sٴL�6��.�rO�pO[�D.�J����-+t]�K�χ�k[ny[�
�߷}#�+RX�C@[�Q��+%�Рy&�
2�8d��и0ʢ���k���Ȁ���k�g��=������������ D����_jIC�all,g�����t8�.M�&+j����1G�8�������- 3j���@�/;7�=s�)~N�6-�5!�)h�e�2*t��%��!pZ٬
�����/�ggo��=�x��/�k��X̴�zܐ�>���m{N�K0�RI�IaN<Q�GxB�W��r�W]sK	�3��G�#�.����oA���G�$�:-x�v�o 9��Te��rb��R�n�
�d��aQZ�ܬ�(�1�/s갼S'hޏ�.T=�g+��8���"?P�r�2$�C�[Oŭe!a�X5&���>c�ﯟ�+�/�p�;��,�?:H�$yN��a�/��T�]:�>�,���\·�'�ͩ>N��?��#c��W.�*Av-�"Zw��r-f�J+�|$���+�0Ƴ����g����� 
#��/�/���.��E���G�i��A���.8;7*ܕ�6|�[J�-:��7����y0{͒�@ >K�/7b�uC�c�d✪�w�6o��L�m�/ �~�K:��.4'i�}.���Ѻt�Vn�S5ΉY��QZ�؟��+��eT���K�+����$7���l������L��I\[@i��. �ʝ��DX�E����p�}��|;k�E͢�G��h[I�\
329��n
���BQ�u7����Y� p�t�@7cz�3Z곱���/߹ �HC�e�������g��w�y���a+ECqDckݜȈ#w8k��hv!gS��t,�v�Um 0x��i&�zt��?.��g�f��%Z�f8�� �s0���Si�3�k⁮��6�$����LQBr���+_�H�[22��6��Ƿ�YǀмЮP���ۉ/�J���7j�{�����T����_����tns��I ����Ι���P
������?�>s��Ü�H�@`m{��V��y�.�q����ݵ�OՃ؏ak��
���G.�o�>��3.jڶ�R�i���R��3'�(�q��?����06��ܭw���_w�@Z�(�Ơ�J�5�-[N��]���9����R+���Y�ݠ�q&w ��׭�q���_�🞣oӈz~��͏�!�]���2�X���n+M�VZ�O+f����m�-']��:&Dq�>�����Gf��L��N%�O�G��< �g[ ��h����) #�����E.�Pu+�*���3<|�Ku)i�����m��Q��Zv6;��{�	��o����֝@�w�F��cu�
�d6?1���WX��]��PM�M�L]�j>S�v%�(D���3v4�s�`� �Yկ ���99Buf�E��i���i���]�h
 ��i)�"Q<]�R����7�|�M�Y�;���C
�Am���zDB�1[��#���z匚�gs�������b@D��BC(K䑍��h�~~�н̝!+ ��[�fĀl����(��#[>���lq�<V��-< ��-Gq+�*&���a�Wmw���P;2?��-��� 7��e�Xg��/6ט	O
m>�����;����X��@ �y����[ ��v�^iJ�kPh�����U]<��K�08V�tm~,m+~I��f������Y:.���R����P�����f��h�WQ�S[��+ Ͷ+$8�v�S��l���%��V�%���ԝ�1!l�m�d3���ȇ�2F9嫶ߦ�5>S�y9?Il�O�%�KX�C�w�3����4x]�V D|����e�Ur���~sN�CBl�ɼt����Ʋ��t��^��B�Xƶ�)�z��K ��� ����Q/�+��S4�w��R[�����b'��,�5mb����W�^��p�A�C�eU�S^0�w�Y���;2e������\��2�6x�_����#�QY����v�����x�`Qq�.�̕��55J�=@�{{���B��'��'ߦ9��I�+ilO�I�'S%?� ��7�S>V�zU ��*��Ƌ�wt��u��$�$��g���J��}}�]�G\���Ñ���O�~Z^�"繨o��;�;C���I�2�+��@�R�8n`�N��Mſ��Ys|�2��t'��5W�M7.^�w�G��Y�eD�A��K��f�>{'�e�8�������g��ϡG~�����\�N/��	��{���v�-r���`a�y�����$k���e��z<�&������;�K;�rv�2��z��=�
�$����7�j
�C��*_�y�>�\�ӆ��$���疕z=�j���}�^ȉ�����3^�\������t^V!>�S/��0m�/�����e��LX� 03pd/]~���(���Pv�ɮ.�����|�9��S��j���]�(�J�{+ES�߀6��i4u�zw�+��^�"j�� ������:����[�:祦�E�z�6�����u���m�]�
 �y�,��Q��=�Ӗ�����R���EL��e�?l�#��{�PK   ���XMe�X&� Ú /   images/3a8749b6-4d34-4b13-9161-5e8eca12477c.pngT{TK�����!hpw	ܝ�\��� !��;���%���{�[���Y��LWUW��Tu���4212B�����-�@�n���7�Un�?�.�����/�g$G��. y7��k��|I�*�����l�l��,��.f&��,��-3N��A�7 �b�G+`ܙ��ӑ��;�dj�$XqE/iL�#�aͣ������zCom��b�"և�寮�)��x̗�^t,�>���ｴ���9�p�����Q��o砞5-��	�G������X����8��	V�Q��	�����t����������>�S���+'nKT��{�ѻ��'��攢���:� ɟ0ໂ��Og^��V��Q��v�m�:�A���<'T6���1ʁ<�	�v-������������|�hI����AVp��༂�U�D�V��u�� �8� [ׄ�*�~�SK�o�Z���I�Lr�vlMn����4j`��R��0j��D]��o�t��`3���ዒ�2�E&��1A�y2R�,���*�I�&9���T9�y�;����s��y|"�9b�ft9�����tD���C���u`�V��s�/=j��0�e!��+�N�ˉq�Q���9"}7��3U�BC��6��J��O� �`���r����6�3t�䁫̴J1Pz`�G?EA�� �+[M%���3i�@E�1S��(Š��������$U����@�rq�,��� "	2��-��/��$d���"��w7eL�~��`�dG�+��YI�?�����S��������b�#&u��]�<%��t��7�\H��3rw��e���/�$<Η$F��C�=�L�/nh;)&#�ƕz��?it紶��-��u�U��J��QS�|9�v��X$*}�����#.[�
���+��s��� �fT}��B��r��g%�a6���y碼�Sl;]?\M.������h�	=t��6:��}~�(�NQAt�Y\J����f|\���a��?N���=0*�^���Sq-.��ٶ1b֎�ZЫ�3"�ͷ��d�)���}�מP�*G�Q&��M4���Bi�n5-��`�������&�x�����_k��*&��O��	ۜ�ߠ�p�=&�5�JȤ��a8���w�5�=�$�� �@h�
��9)$�����ފC�� I&j��)FLx4�[C���o��q�C���M�q��J�����b�����������8-c�� �Wk�
���#�,;����f�0R'!������b�µ��fg:#���4z���ҳ�]�5�\z*kq�����`�]�5;�p�9?�F�=uo�׬����_*|��,/�Ă�Ӭt���#%��@�Vg����\Ҟ�W�ؐ�K���&yRx�)'Ly$@�}��m��X&�5�Y�'v�Ӝ�u>AC�s��ǧ]�sh�h罠{������`sB���R�e'w�&֟O�`1hp�cꮠ��q�Ǟ�⟖�]N]�z���B�?n�zެ��6 ���N0�������d��������a�+�v�0��X"P0�
4�DP�1Ϟ,��7�e+���)��ľD�^w=�t������e�;Z&�i��>��D�Q������T�L?�n�l䜞�>g��M�:�����P�ES�z�M�K�~#v�hH}-���Ҙh>�u�z`fZ�Lu+��A����O
��v�D�,L�S[<M��R��ӝ�}�����a9v��D3Ls�ܒ�(�N�8����g��1:l�p���DZL�����ZSi'����R3�k�]��Y�s39i���3���E��_-K����`HG-����k��dn�E=�\Y��Qg��1��xD���2/�e>H�����Lqx�Խ����^+��1;-�������:�,�kՠ ��U�zsVJT�����M��m��w���֥w�F� ���� �����Qh��>���n�DA4c���-�o���4�'��e>*C��*�w�����K�j[��;QD>'J|�5G2?�ޒV,Ss�v;��+�?K�A8}�(Ib u+:������T�=�b�g�'�os���+��k�M���0�8'�j�<^o�>�m� ShEK�����X�<=��=�oՠ.����"�[Ϊ�R6�Ʃ.>��[޺�a>��/�8#��|�A�0�hC�3����%�i� s§3mJ����u.����v������Ib�OS�
��^GB;vM�͚M��Y:��F�ްJ���扉gݬ��{�	ӕ�r�;��~n��W~Ru���͎;O[, u���.E�7L467��,R��9�&&���g8r7}q�m��z�it�z'���uC�|7(�Wm�B)�FEX���lw�㞔�� 
Z��s�C�V��B?�o!�r&wPlA��nD���Ny]�����1�G�UNk�����rh�醭[�w!���9�息졕���`+W���Η�ۃ�$k�t�\�r.�d#w�B��a�<�NP�.F��՝���l?*k�(�q`-����e�EGo<v���
5X#�<�+k��=�-����ka�T@5&%��雳��z���
�5z��և�8��Ӟ8��Fds�-Kn-N�8�o;��Qa�<��,(�9Pw���Ae��_�����p�>��ݴ���P^~"J��^!��l5��6h=�x���3g1���h�q��F�I��`��j:{퓋����D�y�j�#����uD���t\m��I؀,�nx�UR�H[$ɉEg��� ���Lm��g������bY8�@�=;�i.�v��<��5������&J> t>@�L$+d:*v�&����OH�a��E��;���嫇5fC�]����[���.�ל����	�!.���G����m�	T0��>�a���}�	��/6����Vq2�8��[�0A2%`����C�=�Q�[�Ɋ���~��#^4���	1�� ��	���5��u� ����^_�
?�l�l������5c�9�뤳��"sf�`�t���r��O�16��p~$ݣ������Ƀ�%=��&$������_�mf��"��,Q�%�_Hf���xZ6 �_�`&� ����C1e2;�H�p�F�N;F�������\77&�O���
L��5Jy5��r6�����-�aY�Bf����D�� [��b�U3���, �g>��E�b�#~� �"#-�{옌	N�`�WP��������Y.�$P�tL�--IVf�}�M����;oVc�b ��:���m���VH���(ϛ�UB7��(��rc{�/*$���-��Fq2p�Fѭ9��|D��d
.�R�`�(=����q�t)h<CX<�8��@����%ȝQ~�����1�H��i�d���OL<�H�Y� ���T<���Z�k��,#��`/�4��|���F��p�y�WǗ&��W���"V���a��.��ح^��G���G
�n��g��A6O��%x���4�`�����
�0��V[��6��a!6򏽿4�߸t��Eh=�������2��C��i�>�Y�(G]?x�E7�Y��a �@��O�YW�w� ��ԣ������v��t�a�03���JlȄ�-O#6u��ǌ1����p);Q�Z�-m;��[<x��sT]8?�O\�-�0@��9f�����U�+E������Ck���Cf�z���1A]Pw���ˤ�X������ � �#GC���y�c��\���UL�oL�3�&�&�@���	1�MYm��P䕭�@��S\;' ��S����h��(�O~b/�{v�E�����~EQ��>��ki��z��qc/NN��z3Hm%�7�;������z穣���Z�Ch��0ٰۈ��-.�]��1l���x��]������/�I�7g�����|�A�J[;���Yd޹��:�9Piы�󑏨,|��!�_��w� � ��������)y3L��V>�7�l�)��'��y=A�R��.R4{$�
�kOhO�n=xTq�#��ʝ��h�+]��)K��X�e���#E��@��V��/�Ͳ�X��"0�k�.�t_6�X�Lu���tFF�x�2d�T�����h�@�>ޒ&��f�`!�����8XV��"�:���\�:��$X�^�E��VSU�=��H���<0sbE����\��@�T��������f�;⸚M	��6���<J��:�
#kmؚ
�_Y�
�ue�����yd?{V7/��J�`��~��\��Z)���2���h�hUB'*��"�^�-��=.Tl�ky$��Ns9bicJ���U�z׼.	��^���h��F	�6ö�8ժM�߉��\���|6I� �Yi ���Gb�L�r[�}��T���&�H�|�Wg2��|B)!E�Xҝ�k���8&OK������sq��H��Ts̽Y�J9u����x ]cj�0���0ۼ�ߗ�F�4�Z(~��uu5���[7�����V���%3ѻf?��<�f���@MM�>��^�+�k�T�v�?�VX6,�� Lh����o28�E�(m� �o�P��m5Ƣ9��	��G��.��=������ب��f�*f����4� ��	����4�R�ٰ2A��i2�T*�"�E�)H\l8�O9�8��"T��N*uS���*��2��5pp��7ེ���OH�S��{�c�bi��Mb:��������W�w�d���:����u]-�a����rN��]=SZ�%i�@���`r��(�8�3*��f���O#D��ֶ�u}\����<���!�3Vad�1�$�ѱ��f8�7컹hw�b�^�Z��虻,�	���M���R�i"}Pab��NZ�gJ��&䧳��z �@�E�3�5�p�mȅf�ԼK���]1x,���ij6���i�=�3�Q��"�������b�H�?ߴ�y��ȷ�?a-X<<���@~w���L��=O�(!�/�Mǣd�9�=��:��n�"dE��C}?�vc�FMw��xNP�xz#��*K��������a�ͮ���mn��b��:d�$�
<5��������06Ѣ��	RV\jD�"b/hS:��;��3iᖸf$D��ƶ�E��7*�A9p-�%o|�G����GW>����w�TƇ޴^,l"�IWw6���o#�kC���{�����U�}k�������߯��;x���Y1��n\��"��������(+i�(c��Y�=^x���V�N��	��}Y��Q��c�YV�3�-�s�Ÿ��=�5��a�*��S\�-_Xu8!����tՏ����/V	3 �|����$�b�6T�6?��F�yt؁��L��[�/�uTsy��߰�n{g2�T���l��̲h����A��V�I�V��B�
�?�@�����5�����3F�3���!�*�H�:�-��w\�$t��&a���;��G��J!8����2�̬�@Ɨ��OՍ��m7+Xw��@�0��d;;�kN�4H��z�����
)�l~4O��L�'�/��;j�I{�6H�uh+�$%�{h*%��>�� X�Ī��6������m��^�z↑�ř����P^Z���lz���Mk���E6�zB�%����S��y���U~O�@Y��Z"� �4��w�_�8�}�P)�ױWt�Ϗ��f�w<�M�_iL���$�;H0|E�~����)U���R��yV\\��֐6��8޹���k��̄@�����7�~e�������o�1ۈ^,�!J{���*�3�a�T>xo�RǦ�/a���l�s�4�.���Q�։�W2�$�e7��}�Ū�l�u��Etxi���0�ց$hS����7�����D�;-�'j|ڧ�nx� �?	���"�*ծ�U#y<?Ru���U��j��R!��JC���ad���W�<��4!��"0V�Ñ�����bԘ�f��@�$ύ*Hf�-�ټ�0���,]���E�����Tg�S�:o]HK}&lq!e��&á/2sU"�vI�4cg�܅�zͥ$�AO��Na�y��ę�<u��W��xJ�7������X�rf��T�1�Ƣ��j̘�%�NU�Վ��b�S�j�v���'(:U�����8�&�Y���_�H ���j��;uobv��;��뵔r2����`�t�;A�@�A�)�ʸ�]	�h�篊{s�!��
R����}q*82!e`�# �"^��2*Ppk��������QSM����T�_p@�6%*��i��z��8[�(�7gB�?y
���"ѻ�"s;���gĿ�9q[�s��C?~���Q�)ӊ��e�7����׎~!�X�
�W�x�r|�r�4NJ6~f���6��	w�uݫwU���y��&��AqMQ���y6szAt˷/,>�s*#��Q$ ��5"{� �(��!;�n��.!��.j���wq� F�G����Z��T`ո=�CV�H���"UYkw=C�����^�l-C=ݞ7�sQ�?z��]�΅+��r����WQ�
��s>�͆��v9[�-L`��i�e_��0w��6�����}��j�O�T��e,��w@f#�?�I��C�1V�)W�zO�wh���r��R��x-�Z�D�>�X;kRx�U�O�{�_ӌ(%����k���G��	�xN�zh6v�5K��u+�v^1X�ϑJ��S@2�<B��f�T[�]v��L�U_��`��!����.��%3��@(���=i}���2�ތ_a�_#� �w��v�07��9����,t��ӌ(;�,KT����츈��V�^�ϔ��ϒ/���]:#���ƃ�Ơv�0�a��V�%��ՍȻ��a,�p�J�~N��d4Q��y�zS7��8^�y�Jsr+4k�<�߂�O���0��Q���Y�5�9�5|�c��|U�XA��0gm�ݡ��d �#����q&�O	.S[����Q���!.&�ܴ�NB���_�l:�싸�ͬ*�!5CW8�L�&��M��c�+�V>`,+��6�-w.iT?ۥ�㡵KM����^�PK��A�ע�$%�ƷRR��V\=�ǿ�f�ͻ��x���[�qjW�#0���*���~D'��x����>�X��W p�iy�I���3i��+Cײ�y*��@��嵟7
�g�bEj�!�|áY��/q[�ו�~��⧂vۥ��l��K�,�19���û�n��Wc����̷��r�#��Ǝ�sfҩ�����2fԫ�����x$eTk�G�S���"7�ψ�[!{>�JH��]s��_Ⲻ�F���AV�_�pq�n"{�3K�a� ��2�A����\�a����lP�[�|´���Ba��Z���@����?�H`:�S��~� �V3N�~ZcD�/C�՗:�OL�q�Lfy�k\e"%X�sd�P���,]/�#�䡏����8�R�YGD��
�&���eh�Zy����Јc��H~*�ǊO��<����u�Xv�hl��{�d�7�Z'�z��/x��c�P@��0�4���z{���J�8v�ѩM�p��E, 7�Z�(��v?�6r}d-T�c�[3%s:J�T���l�8�d7�o��0Cؔ��u��*#�E;6)��� ��b��-�f�I�o��
ε�O�������{A\���%I�0��k��%4:bf�)r����W3��)��F5~���}������T5T�$��荡����b6�S ���q,ތ�D��I��"��f؎7EwƊ�@��:����;�i2W"�n����F;J�G���i�` v����z�D>��钡T�7e�"��ܥ6��m��E��q�"���R�/T��fc�<\¯��'Zl�a>h����2��VRKn��ʥ/zޝ3�Y���[E�z�H����kq��\c�s��VT��ޓ�f2 s��{�$Ht����=�ċ3iE��؏���k�/�V��v����j�̠^����H��#�˴�PY�����Jlqƨ��"̂�\ݔ~U�ʤ��x)��=�8������a�6�F�=��M:�3�uZ���g`��E��SxZ��@�R��'� Уsi��=���
�n�Ýn���3�g����ˤϼ�]��^�"v|�H�w�8$�e&�&���ޅV*���?%��W���o��o���6G��9����p.b@�����Ⱦ��z�]t��}�V{S��� {�q�8�\�[��q�U�C� &ݭ� ��6Z���4"����u�%�3��T���6�+���י���a���ڕ{��f�g����+J� �R�L
R��Tr��xu��O*����US��[�N�;r4�cy���="��䛗��t!���.�/��^m�G���_�P ��i����^�۷Vk�:������e��}E��q�m�~��K�q�KŶ�^��G/BH	�T5Ԉ�"�߷������G"��؈�WBD���@m�\Q*D��\����|�����9�ɧ���v���[��a\�V��D�l#�([�հ��H �5ta��ב�~�+�#f#\�En�N���!��`.=�����[�*bk���� �K�s�{�.؆���)�5�� '�n����E�V�?Wk+q���N[�I������R��l3�	ե���9�h����c2B�*1�!��6�{-��U���6�i���<�m�0f��9$1�J�6i��_U��~�
��;�͊߈��|���WM$f��ͱ�v6*6�����j��]�Gh�X��d��[��{e���L/�g���%ŗ��5��H��jhy�=U~���A�@��~�\�g��W��S�-е�"�Ht�M����o�lqM�DW��P���;���$���c����+�Z�\�oR_3��ΝgꏟUic�mg�N�J"�b��Zw��n�aDt0��6���?�"	����X��Q纏0���7��!���ژ���b��rb�sƝ��vy�F����F��*{ U�� ��/�%�C2ѳy%�C������&����+��	ƣ�l��%e�w���q��[w�6�fpN\>�҆���0�pa����5�93�5�����5`mT�7�%��k�e't����V&�)S.����P�>� �7i��T�DE٥J�wu�A��b�bi���JjMp��@'��K�{������M6�w^����6�w��B��������<1�[}��a7Ϧ=��c=�^��k���9�.`h�u���*�A����Ogf6m�2��Tm�M���%܉�<ڨֹ�#�����^mPs9	�;ĳ�ֲ,]�w�����ؓK,�Ϣ���u���yZ�}��sNA�z��2S5��F0+�%bX��D+�r���L>�xx#�|L�f� ���
;�%P�\��?��D ��F.M8��-#(�}�����f۽Q��>{Q!Q��(&
�PW:}�ko��f*���7=������E 7��?�ObJ'z�)�|����1��S���_�o2�c�F�H����n���%�Z%�J��+c�X14��C��I,���J]�f#�uZ�A�O�b�c2c�|���9z߲�o�w��$��Z����9W���Ut�揎x���P�ы-�W3W��uR���Ⴂ��n��)����b��4X⺳Y����Y=�u����4/Hfi�Ko6\f�cgřM��v!r%�ɉ 7��̛��P#gy��B��1e��3A�v�k��
����ܻZ�F�.n�϶�!����V���q�D��{����كb0d�Q���s����|��t�a�=}e���o]u{��0�z?������o�*g�k�-�T�*Ǿ>��s�
�(��|N����97�nC��vE�XT�[�@EA����%�oe5j0��f꽡�RJ��+���|����������~�A$~�h9�V��I��L|�{�5g?���{���mL�W���K[>t��sE����&w)d��iλ��P��#��x�5H
T4�[i��'o���n�ݛ�x�!�LF��C�,�3�x9��z��v��S������Y!A�#��@b��_3ŻjH����G��yj��m��R�_8��|f���t��x���7W�&Uh"�L�1Ao�y�'p�L�]b��~N4`�LN��I3`:>u�>n��򤠷!�cR�����
HD�{l���VNfcy�n�[y�|�EG��(�ܖе7O�`����_�b���"��|B���q�q��P?�Q��_�p9��m0��j���,5�M<�ϋ���%�a
��o��A@T��d:�C�	�]�_�n�nľ�s�]SE�!��`p�%�N��X� d���((���9��-�_h7� >9��ϣ�1r�>�F�.��|ۊFi�:|���*+�YFU�pa~����2E�a�T�e�#��%B�^M5������L˞~϶��cr� 7x�X;*�����qj+��'#��]vТ�ϕV��h�U/�O���r:�K����	�YiJ�!G�x��i9�ې������&���'�����r��]��?r�0J�2�5pf�:f]��g��ZQ�������eX}��D�.�h����,,�?݆��?�af�''E��	����U[�d����m��f1�x��\���.ؿ����Cqq�F���+`�%Ĭ�6zd຿:ej5_���Ɲ~���lU�}��X���$��WK߳j"Y)º��9�Y���iZ��r�ݘo�����ةW��	� "�jd҉�*����fL�jθ~���_2�ed�SA����6�CB�Ex�t��ˋ��©�嗫��/"���U-1@g����&�"�ˤ$�Kfr_�țk: �BU��1���ĸڳV&{����NZh���Nۭ��&*䏦/����f�տ�I-]�Z?�`��++i�sO�~�O���L3��M�6�Z��J݊�Fn��d�8B2��U��!(�j��V����%D��.냣�1���tcW�l�U�6��H�m�N��A�eۗ��ni'�M8�DM8�&7����Ƭ}$�^;�m}���4�BW8� \ԡ@�
C�ѹ�� A�P��x�l,X���!�k����D��l��R�O��ΰSH#�b�?�oV��߉�V�`��B��`*<�8E<�>?8M��=l�9��^�-Y��s�N>8�6%:��쪏��Z��$T�~L�v|�}�_��f����Z��s�1I�_���e������9e���ɋã{իU��ػ�L7�J�K�Fú�(����7���&b��*fV8p���4<�S�N�{7q~���9=ao�������������54�'U����!Ͽ"��H�+�P���L"�.a�m�d-��L|lA:�;HǺx�p��A[�d�Q���[kI�?�Ӱ��:������	�R�-@�{�C�H�p���ߑ���$�f?�ә�����h_�h��˾�Q5��FZ�d�n,{	�lH�H�m0�tY��S��DZ�d�� e'��'z���Kv�}��*���'�8���9�	��1�HS�$�\�{�*`l�;)R��'''�]HU4���������߇���K��V�;�	p�F^a��Ǟ����N��o��4�S��%�s��Z�>A��ܶ�L9��[wEZ	ٙ6y� ��M_OO�T�`/=� ���,�p˕�����+�i'l҄�p%o1�Z?n�2z��
M�pC[���^���C�����G"�Jȡ��;�>V�"��'��;%|�Q�$f@�����edd��l��II�hl���Yd+���D@1�m�9����O������W<r�I�Yj���S������aG����`���a˔!��厽�G8[y�:ֆU�X����\��:TV<�����}X�=,�D��[͝p��rpmeDM6w}kr΢?e��n�W���mh�7�,7�s�vns2�y>ղ/#�ޱ��3$����-c�xP
�C�G�3²$S�MM���w<s�TZU%��Ρ-Fr^R�H��b�P9K�a��:�XߏHk�Xd�ux��^T�ܳu�8QkB��ޓ�Ň>33ST�n�GE^�����:ѡ�[.wx�>N�<l�g��S�\C�����:^/�#�)��0H��b��dx桺��?�[Z��T�?tKg�2�f�v56*�c|�};\S�d�}f,D��9&w�#��
*�*,U5�<�W���$|�GW����y�P�>U�BLdס�DSs���U+���Y����D�zz�%%��n
��M���AKdD�y�?�Vhy�}��t(��������ҷ�p	�DDDʎce�z��m|Zz�*ot���ο�n�-���A���$	��mr!����X��4�����e���И�>��,I�
�T��·�����S�b)>7O�B�V�����y�s�k��H��7�T��<�f�Ty�����#צ<���gl�떣�>a����Xq���<E�w�{�9p�a���bB� V����,Gcj���i��C�A��{�đ�J-+t �N���O�I��&V��њ��zbti�'��7�o{ٺ;S2s{���Ą��n?���'��z-H�Kg���+��o	_��-�*flL�NoQnZ����3G[��M�Ύ9������?X)T<��Ƀ�j޻t�w�o���>��36p��8Pq�2���ٺ,��]�z(\��	�1���Xb�[s��]	��>�p�c��H�i1�V?*i�޵Ӄ�X��Y�3��n�g6�'�0m}<9QaZWb����A�
Ra|j2Ua���j�T�*El�9�<q�ޘ����#%���a�̮u.�F�m�j� �	��qEZ8I���p�]�DZ-�֮IHK0��k#���$��p�4ZíI�@�"8�f8_�	�[_��&��D�+4���ՎZ�wF��,�# t�A�r�6\�M�LJ�GNB�R�{�z2���:������y�/����|��D�%M��u���\A��('�����e�M�riҪV�E1��)��}-���S�Qn�
9L�֝���<�6\�%N�=��1��E�dbŊ��A.��`NhM@E$��}i0U�BѤ�䶹�A�]��铂�B+�m,!�^��O���NZ�9Y%��e��Z�������h�ݛ���ޡ$K\Mo��N�[��xz�;1ҟ�p�Pn�*U��>;��b���E���^ƕ vx�!���&�Q����J&���9��4�X�Y�?I/7?�h�~��S��D;<y\�c����rńAYU���Ђqώ�!J�X�wk$Q��6�J?��qT Q��
}��~�~�wo�*0��7��@���0^K��4&	;6��t%`���:u0��#��X���O
W�a�1(s��T�A��4(5��ԢϢ��-Q���h['�@Y�?6|������U����4m-ָ�mX�>����k��4H�F�jG���.'���v�$����d���L��H�0���2��_q���L�_� ��������w�U�r�
�.���Z�0�G�-%���ʒ��aV	
�<�̡T���7���Z0�X�@	�0_͊���se rN���n�R*�Չ�HJ*�Wuq��������a�.a�U�`����ס�+g}a>�ytX����P����P]y�	H�{D�����WsV�`�&���e��IFM�:0�d������b&���I����c�<��y�:~b��`�{cZ�P���0aP�m����o`@�f���`#"���R
�_��0��$���gk<��c��OR/���h�o%c��dK�1BMJ�8�7��X�Cv��0i�_�8<�=R��*r���명<���輸ƻ*�E_UF�3�k~x���Qc��z9����]��o\SL�~T�p8R,�#�a0:\;��5������m��x��$4�v�2Fˋ����B��W�M}j���7��6�rm�۪��vȦ|4!�v����c��=��{�xZW������Bl�=`	,v�dK%}�K+$����ɴE���v(4U�u� }���4�g�Ž�"�Xo��a���P���9j�M؉Z���;qp�;��ʎg������ߞ����=�@�f��&P�-� il��#�u5�?F�f�ʆX]|��3j�\ ��jx��]
�J�
>�}�����ZI��@�b��@��"I4{���z&�@�'�%O�з:�2R��ҏ�7�����>�R���"d�ڭm8��n�L�+�7�������wg�Q�Q��w#IF(uw��ɚ�6?�7�D>�R:��3>o��ǝ��-�i�N�َ'�nK �����s$��(b��#w�qv°c��� ]�O)�m�P��E���w��Z��A�yrʖ?�^ġ����&����Wx��%77��_"$�g1��-2��	�=��ݝ��tb_�Y7$�E|ж�ѧ�P�n�r~u�S3�ޅ4���c{{q��l"�}�������"�Uz��Tħ�?�D��٠"��-��� h��,����^ �����׵ߘ�����EDD�O����-Ėe�oݠ��'�k������[�qp�X�266��%P96��w�������ʁ
 �5*6�=��x��*�D*�����>|������J�Ɖ��SG�ViB��	����6��X2���:d�_�b��i;~���^y�~8���)�5<�l�_���������}eT�V��pm<e��V�Ձs�|�_&�qp6�ئ�	!����Pn��38��GQ9�9 ��|ݒ>�� u�u�I�|�����Q�W�Qe5�����l�DV7ˆ�Y_��5�38��Qj�8�Ng�����Z����М=.i5�,W�_N����=��w�`�S��j�w�W,�����M�v;л�]´t�zyoo�����އ��;�����T�4s�o�ǖ���&�	Z��`Ѧ����&|a����)�M�t���F~HU���_�Z�����7��((KO:�K1���v+-x�/wTZe:Pq���N���Ԃ�'�?�~E`�|�,/W�r7�S������}�g�����q�^�O�ꤓfñ�4�l���u���c%��߹�,G̔jo��v��T�p���$��&�_����ٙkD˧��>��,X-����=w��43�7��ɿ���˓����i�-i��S������U��A���MXq�@)áyyoq��r�V6����Q��T�?.�bZ^�Hf({��'�:�Wn��d���/@��.��{1������Z�82�[ݠ�2׷O`�e���0���d���xxp��h�Kd��7G0�T77M��̄^/�X��De�-F~m$��N�:X?;%}���3�_e����{����u���y�W���W�?6j��MDw�6z���	�!�
�#����;���>C��Ԋ�0����}�`$��}��,�"�N��)��}a�'c��U&��e``@��d�2J�d(�c)��Bʠ_~��$�bF�,�����G��Ɣ��K�������ZR�WTݸ��$�_����.���h�>���ml��ztW�z@��a&�O,�{���۾oC�ԷO�>���/����u����[h�U䧗�*���==��*%�3���p��yv�C-¯�\u,��ur�wha���^TWa�vw��M}wV:�I���+R���|^mϧq��7�R���m�7F��ӌh�Z'�U��f�qF5�"��͏���V���！8���(|��?`��?IZKJJR�[��͒]�>�sEF)���c=?Ҿ�仐��b��KB�����k"*J�%��HτڎX���nD
E	�[��j����@�����5�f����/zǋ�gI���?��g	8���������61�����8�E1�	�QV�|��QÂ���<@�� �l��;5�����)~���l�~���D:G�K��a������e�}���%#4t�7��0 �4IG8B�Yx�p5���?U,q�(�v��t������{`6qwUd `:c-sT��3>b��o-]�$N�@��|p�3͗�*��gc,�^�≸j���{	Q4���y6���#�]6���)\��s7�r�����0��0�b 1 555����@&��>��7����ї���R/��0]�b
����2�{XC�K���e"�`t����7�j�Ł�Kjĸ0{�U:����� _ҭ�~��6�
�U���"�O3a���d�ݝ�ra��{l�,�HL0?W_U+�'�.++�NA��1uz�=Wf#j�\�c��yB�i�u돂����I��%O��fZ@͕efXy-�

�G���lU:L_""{7޻�r�4Sz%�-��E�Dc�q��
�㭕�,��k��ŷ}���dmxR�!������_o������֔j��7&�-��b�(@�����-�%��c7��~��
�Yl�F[�+Nz�*��b3��-qe�5̑��"����8����:򅴿�P��ob 8�/g���0�Kq�	��['$%QPB+����[����r���\��a�)��j+���	Z��<�׷&FѰ⧜��	G�.b�LMMa)*�flĖl?SX���0K�u�9�W���sb��f�!>�ԧLT2bl�0)(����Ė�C|`]:?ds^A��ԋ�ɶX�,�l%�ٲ��
R:�ܓ6�2��>��t�4d�e�V-5�>n�
�a ��x��l�JnI	�C�ޙ�R�	a_���Ն���_��GL�E0�M���lǀyS��"�/:����0,�WX~�???σ�|�������Qq4Q�8�� !��.���.����	����]Cpww��]~������������e�ԩ������h[m�Q���	��.{�~T�œ��w�ăv���	��YFj@3Φd���崴�4�k��	�A�JJJȝɪXA@� ���n�N�M3c!�DF��i5�K� 07��m���Y�Z�4��=8%��ee���E�+n!�]�D���>q�A� �K~�R��VD�K��S��0LK�y%�3S�1�^�M)�)>,���1]*��a�����f����u�$#=�T���o���D��R��u��ђ��SR��oW�){�Q�$�2 )o`�v �.�0�:��0��Mà���P�&EO��F��Κ|��|y>�Jfϸcr��S'r��kZkx`��dP���u}ĸ ��o���t�� *�Jgͱ"��>H~�qѤ �x��|#�����:W���'���aR��aj�/@~�%�C'd��^�/�[A{T3l�ƿ�nL�=�\B.Հ�y�����d�A��w�ݝ7����nD�#,�2�J�A���N�Oqm��~@�Q'�>�2(I*E��(;�7T-�A���]&��&��g�� ���������w3k�e�y�fff��C��������r?yb�����8�w���R��~�m��I��F��%.��-��;�oIo�I��|@h�-�) "P�%B.%=���W\�i��O�vm��s�0`�FT�\A���@%m���#y�XN��3ϫ��A),0dw��n6�.�3]�l~�_E2�]�P�x�:p+\���$�Vt1�XAn��^��e�!V{.L��	�
�n
���j�>���s8�
��0h`>�rZ���!����OB�z� ���p�"|@�8��1��r�<�5�3�[Q��A.��iDsK�P�cԤ�[𫻳%��пgŤS���!=�JI!D�-��ss� C111�",�w44`����z�$���m�@�KY�Q��W��)M���M�?���(a��7ݕǓ�(}'���k�LLU�������

���|i�uV����;잵��l�/�` ���E��Q�����=���\��Ny�������w�4 RjTs�Ӎ0]�^��Q֐���Y��� �=0�/��"^���n��JJd˹)��4���V3e�60-v�P@����<���_� �=��]�~�6�B���[cy�p�p�:Ǚ������٩�Ed�]���~g��٧1R�.�*�$%c�ۃr�]�XXP��C\�l`�'u��j��Fkzu���wƤ-� ��R���|��w֓��#�1g�@H�ڹ.zE 1�#��ń���d��G#�e���"S�2�ܦ�?��5��1�T��n_�!U<S�!EBN��/�=�@k%z��\͍�����Ϊ�|�s?"5����)�l���L���IYP���<���+�2{#���뷞��:�̦#;pj[�9m���UP7��Dn[Z�A����<k�d����S&oo(�� �2��q��F���vz�tP)Gv���&�x}|��1~V��[����z��^�@~���6#���@ç�F6�":᧧u��6����e��)r�˘UCcm��Np�m�˗�:��Γ���
>j)�� o���Gcې5��C+�9-T2y�54�`�O���/K��S/��_��\�Α
5���P�x4mBǠ\V?��:jL��լ3Oc�p9mM��,���h�'8��`��%��*l	Y�����	a����o�j�{��$�.�oE�@	�C��bH�^0�K,�9��x�+c��y=N���l���3��d��.SV��O�rrHڠ�[6�
�zu>���n],g!tׁ�U�A�������L`DX��sr���iݏkS�U����	�㞌i)"DId���f�ٸ3�l����O?��*�>�����=����unT�����W(?��+6}�{oC%'WA�+��h�(���f��3���x��b����B��I�D;j�wӡ�T�۾nj��qFDZ}N� ���*@N�2rb+"��g�4<�늩���
�֤�G%iW�J�+�#w���L@7�=^��]�w�&7��|�Ә�A�mw��l�L�<�G<��y��'�M^�e�Ne#�SU���d�*�XP��ْ�g��ӣ����?~���|H�����߭���|d���#�Q���~v��kOa��uْ��y�)�|U�+�~2���3DT{~B(W]�[�F���w=��Jr�c�X�-p+���_��y;��|�C�?ؠȍ�V�ޭӜ��%�}Ųـ� 9%�٢[@�܊�&��E�'[C�@�c$���#n��DP/Z�R�Q���/��J7���׼~ϝ���\��v}���	���n�hmm��r_�"�c� �ux'{!��J�D��(H9n7�!��D�e�D:,�ȍ�����o��
e�T&T,Ylr�bm`�^޲ �=]�9�5WB^�>�v����d�egl�?�%��}xX��.�H���ZE�%�$��m�UU�3Gl�	F����#�.3U8�`��\]�]�
2���jŮ�&��wS�����dڞŒ���&�da��B�/�=G��4��������IŽ����.�x�W+u?�M�p0	Ą4¥���Ƣ�����Ѷ�<�w��f�|��$��
O�wf���&�6� �+A8Юȷa(��F��c���g�@���O� �����h������6ok�C��[���|��5ݱ-�����D���]μ�w�C���%Jv�}
�P?��;:������µ�q�V�y�y��<����/�ǧ�gB��� a�\J4����1wG6�s�KL%��_܂�p�F�ׁ�Aĩ@��sH �L���ZG�L�r�"�(�?I����`��cݲI�%�ީ�����4��s��ʡ]~C¤NJ~9�(G�[>�H������o��e �壣b���[�@��:y��ڨ�|}�p@�	>Яs������O���'6�z�u���ۺn��[��q��M�&��[cs9�}] CuN,Q���=`��>R�ky�'�hnfn'?������L���x���3�e��� A�kx��vU��\�}����n��q�̉WE����@����?MMM���EKRR҉#���H=�%�#��������C�~9�߫�)���v]�ke=M���lc�v��J55���a�rO�8�K��Ԡ�p�/��ߊ��oW�c�j��'ĔS[_�v�ҏ��e�e)�ם̳^���/��6�ո��\�����G}ߴ�|]�&�] �����I����ٯ5�ﰎxQ��e+X6�9�7O�J�v&T57�Y������H�4��1{\�~0���h�,�G�����w��8�$1�����dT���#���)����\?t2��6r���M�i|!GL6~��[
5�"��N���!Xk�W���on��>2�g=���a�1we0	Z\��������~�ɾ��*)�Ĕϟ�d����>$�kr�|{~������$������{i�g7]��
��Z)�����+_�� P�fcǐy�Ox���;�
�p=�OgV
Uϸ�~�et�g<YM�pw��z�N-f#im���7�=o���V>e���L"F:��P�� 	p)�#��N+�!Bzf1������m��C�J8�8�������W.��f�/.
:��;�\��'_���A�{V�E�����j�8+I�y/�5m�bgi���0�����*��U���k��3���� eq�{�~��Y^|+SÞ�q���RɈ�\���y����TYJ,z��~�G@�I%�d����c+�"��!e�9�2���l���cM�H9C��y�4}T��ZH͏-"���yh�O���ikr���9tJe����a�%�}����uVo���-�m�f+1��	33���Raf?�Nܫ+�S�ff��|d�V������Gvﺼ/e~[Kݽ�}7D���d(�~
е%��Z2�I!v�|�"$k>�~��͉A1JuT͈� �N^�Q4��n������ƶ�����(i-�����{�Q�H�Xs�B3�"�O�P����X�M~u�;s�����L�x~�O���P����I���+����JќQ&�عeF!��t��p)+�u�9w{�������e_{-`�%w]�=�ҭ�����Ff�|�*��,<='wt=�:��,|�q��w��x�@'��e���ݱ|JV�Я��c�q���	�S����%��@�RҰ�����\�2����y�� ���*��/V�^U"@	���H�'͔+O�PW�ՖY/�f�.���D��^B��CTyg~���-3�0�7�˴�K�M�u��B��P�ϰ�څc��z>��{��B� �/�
ʫ=J���9�@�K߶��TX�i����y���i��;�}�ͣ�fSֿe ��\��ݟ�I�>���R�0%$��U�{���Z�:.�� Ou�-�zos[�L�W��n d�.^E�x��X8VX��f�N��򓾈8�{bz���z�߈*Tg]E�;�ZUZ|�VR�+QR/�Y{R�4���߭�G'
~�H���Ur�h+O��*����!�OjB~�x&���]u�2��N!���'���D���2c2;�9�!�Z�~|�B����5����g��i�!���d��=�����d&���-,`J�>��#Z�Xv,r�@��r��K�[����{��L���EUcK����O��D9L}��L�q�
�|������q~�$M���H��_���5�W��R��ӱD��HnW>XCߖ��0hǏ&D�?*�4/<���kn�|>Ka����H�.�/,���!�C����K��`�s�+��E���<S���>4����L~�}�~���n8��r�T���^h�f����*�C��aܧ�*�WFf3ˁ�Q3�~Y�_Dv��@'/����_$�s��%(���XK�e�E0���6^�{�1n�w����>�kC��k(1����X�~��{���$�0�3��b��i�wR�����_��:�j�Ca̕��|dJ��5�o��V%�*�r�n��y[���j�����fR�c�/�6>h�c-��7�-�� �$(�J��D�!���@o���~�>Q�����b0��y�+t�u�l�@��6p�U*���D6>�МL����h���4}Cg5iLߍ0��1���|��H&?����#6Xe�7W�AR��V�����&ȩ��lㅴ�� 	a�H:��8(��0P鞍MN{9�L�׍e�u��YT(�������^��%;�{R�t6�؃:�~����e��'�(=+�W�YLda��bz˶�S�� Re�q<�6�i�j� ��,�U��V��D��Zo�4��/�W,�r�`:�~Zv'�.���c1���Wb B	S�7�O=�<	�w��>�� Wg�X-nO�zN��\�����&����654d�����!#��OM�� ِ�l��W�tuNqԭ7�`I������{�4�j٤�\�D�/4�ߞ�����%FEka����5z���T�����N��ˍ���7���r��G'�MW)�i�޻��C��s��;��&�y4U�#ݼ���E��CRN��I��鞄X�^�0`����W%q=�ͳ��-o����4����������o�?Ax�TNit�D �X6��P|�_	f�à�:�s1���C����
t��FZ4y�����6��3qw�m6���ٲ�#��B�CN}���0�ٰ�d����E���O�˝�mO��jK�z�0� ������������� }�5���:I�#wrnk�\5c�lC��	�v���CX�����v�Lc���ֺY�fD9�;�ŴŦ2��_J	t�9�˛h�afk̶�i�����]
R7[�2��L<�	��C�A�)�����/�I6%ByʌTt�c&c�?�Z�U��>X�g���"#����J
��� ������+�_�Y�j߁���Y��sx��Me�l�7`ס�E��p�\���0�*>�4��"���?[7QKW}��NռR\�Z� ��\�B�	^�dO�3�e�1�z�� �([����]�s�#>��Y�_�y,�^:La�WyI.��l��֣��+G��{�lG֓'d����֨V�a�+�L��&]� �[qJ+w?[=]y^���U�N����z݈�VJy/��՟ѿJp�3�6"@j�뺑ٵtxX!�\[[���p��8�Ƅ�|%QM�k
.�<���àD�����|Eom�,�x��I� 3}ϲ���L���������/1F⩮�1��B''�N���#�jhI������U����2�8@l4�'$�n��c�^��h�՝ɦ��B�K���$��������e�5�d�e(H�CxƤ�A �1U�JJO��]�M��x{��W,ώ������ �������B�_i+��n�9�t�lVb�O+P]_oB�Pﰽ87�f��Q��L3�̌I��+]���閣�Z�0��%n��V93���*���{���p�	�G3";L�Q&��3o����ʪ(��o����|ؗ��O�+�>�56"N���l��93�$ʦWܦqgX���GGaU�Y[\��=�ɤ!����Z6E�W����\��"e����R���6���#N�-�l��l�Oy�+;y{�����W
����}@�h
p�:��������9#�����8�OI����zD�/�p�$�����{�	�"6�:\�P��!��{7�s6�	�m��~5�n��׎�/�~���tPo1��Dcj�O��`�q�H-�"�JⅼV�ۆm�{-�E�U=V9����Y�bj�a`�8K���ۉ���If%���`��`�B#�?ӴbJ������ �|�1����7���fj�&���2>��G�6�H~V�5ƀ�x��*�[��vY�R�	����H�!�����?'�̘�JLݦ�����Nb�N�|�}/M֚	��O��tϐ����Dk)�u����_��)�	���L受�D����*:�rU��'�⽫���YA����!�������>{rr)�oi�x�I��2��i����o �$##L%��y2�%.夾d��1�h��<���W���`q�ц�a\�V�$6;`�-�� �F�r���e�uq�늎���=΂��d��!��ڂ1཮<
����3;��;���<���R��㜭i�������/ �9�1Ac��;�2_/%g!��0�cx>iNGj`��W3ϯ���@�Zmo�������w�������؇3 @�;5�ܽ���I =���~2�d*_N�/J�s��p~��x��n#�J�K��34�{/���58A8�{�f�O��g�ش�C���ۿ�f����/N�c2��Iu��i׾Z��e߄�K)�;�$�E!��;�D`_��S��Fs�G�� �vm�ˊϪ��c����)��z3��ɑQ��Q��G��
ڂI�arE����6���-��߈�n����2������3��R��5C (<J��n����#�(�|\�7�'k��Sq<*{���b�D�07�S�!�}��)y�E���;;����7��2���h�P���SCEG2�G���iLP��4��	O'���gYO��V���[[����>�/q=J*"|�oL'�N��ɠ?��8�C�r���O��Ɖ�u�+��d��������[�{4��a�h}�Jb� ��n�$�~H��ђ��6��-Ւ�rD��ಚ��x�܃?�5�y;Mx��VT:h���Z�@�4����D,�n�I�Ckpd��>gcN�L�rVuW.����?�kԎ�9��~� �:�6��4�l��9м>�N �&X�2c{qrӶ��Z�F����3�u�]��XO�[Z�+�6U5��n;�#A����`�(V�b�n�2�8��ܳ�/�,;'�Y�H��i����F��*-=Ъh]��s��姆��x�5�H�>���n�����͟[��A��(�E��Q8 ~��߼J�uG1[�<m���C��4���<_Nu��5�m�:NM���2�t��iJ�� <E����#y-DUV�}Wܦ�2�j���ݠ}�^�̘lh���`�g�G��NB��<��66V3w}*阦k�O���=�w�lZa�p���Y�����k�>DZ��O���sa��]��T Y�n<$��+]�g����`Gj&ԟ�g��cڪb�e�=��F��������}����8TWͷ|z�����`P��������C#Y��1�&�
�B�ު�m�d;ꡟ���������4nY�gAO�D��C���g���.'��Z66�I;��m��f�LV%�n7���+QWhژ�޳2�Y�g_c�3�L���p_	;��d��D	�
�n2Ԧ[�h�>��M|������ąʘ|D�s����O���A6�zm6ƃ�zx�Ǒx��Yv_�2
������Se���&Bڥx5"Q�d�̃	�R�n�Kڑe�a�a	Nu�
��p��pͨ��DeVf�� Ŗ���kCʼ��A�[��N�o�ї�5��Q-��K2�ق>�vc�Y�z����i�����2�#q���� 0�ؽi��$�˻�<�tý�h�;o/h��}�1K��4z~��i�*�}�Q3u�d�}�c�i�a���Yi~�#,�����i4Wg�����_�mFT% �Asu�zh3�k�aKKwd�F��|J�8\�7[�f���|Fy5E�Y�t��_y�6��w��J)h���
�]�b���&��˨��P���c����)X�	�V#�����~�̩����>TBLGu_��0�R�OmC��J��,T���y������0"�j�MY�U�������d���.��]���oR�����oB�����!ڈ����m4Cl���'��N�G�v$�3Z����J��PݩGg��5ե?Jq�8+%��v���k��U@��Ȋ���U6�S4O�x�@Ý�Y@�qѾیIٿs<̊�]Q �Y\a�9�I|<���]���R��!�g�c�jj�΄��o8=uT�=Sď�2m��A+4
b��m_Rړ�K6�,U#Y�����W�)���[��*�{d\{�3��1��e񙓩�.ar�fp���6!�̉�k`}���h�@M`�չݿƫc��+�;�����=�x���ڦC���©3A˫LV���5y��O���SC�6��o/nd=Zy++��Ddw�4��k��������v3���>�}ĝm7�޸O}Z�d�l^P�.�R���1��PT�Z��n�� �7��\!/r�d�mM��|��G1Wu2$Ku;�Ӕi�4B�x|���h�"���4�O��4%� k��7e(�9S�^V^-9��������_��c���s2�9���ȳ�U]Eupo�]�?�u��R�����٬t8��	��	�y�&�qV��������ὑ
D ��h�ei�(.L���\$uy�n��#g���˲�ɖ��"�۾�YS� <�m��II�T�m�q�c�ߋP��p�l<�jK�_x��cӽb	M��A�~=a��yM@C�-S����-�y�ŬB�c"b�?�i�L���Uvml��}*�qQ���4����;$�SȦփ��B`�5׬����UaQf�C��,(P�|��
��u�a��#�>��� ��D	������U� Sr	����n��h"x�l�u�����%V�`;[�'r��SIp��ȋ���.*�ӂ�n�U��� 2z��K����{~-��ӭ�mT.�����n�C���k�p2�5�*��'8��)I"�m�����N�2R,����Py$�<m�W��Y�>�|j�[_Xx�>�ސF��~7Z��oxg?�<���"�8��.�q���V��7#9���e�M���'����*�A��VP��e�,���C�4�*WW��;��W����A�y�È��[#b*��+��@E��P}�,�h�>���@4�n�_�	^��#�|�#�G�p�wK��>��5����<K��v�z�8t�ƹ]��'q\q��OΎ����*���{���G�-5xjcn��s9R��v�2�7lc�����LH�q�����i�>��i�@w�w,�n�H%P��  7]\�c�v��	����J���n��ߪ��6����;#\J��de��u^ob [Z�,h����C���{�ײ��q^�B݈b�	?SD����{���M%�I�uj�^<��9�ߓ
;��	L�^��G�܀&�ny/����V��ǫS(N�~���FeT����E�*�#�Hr��j�c�^��$ �u�IYt���Z\������Đf���g��������M;j�jS����pn�$*�5����,���0/��MuyY�_�[M�������W9�,� �I��W�o��n���X��ݤT���A/<�KE�;��{+�p�S�3eK�wK��L�4[<���ͳ��n ��}Y���.Sfl6�� �~�+ɪd�yf�,��ݰm1�k�"e�(��C	5?.~���,Z$�@}��3Ķ~���-n�O]���tTY���Y�0t�&�O���S�u�e���Zk}I�b�~rU��9}���&/����>� ya���XKU;������{o������%ѣ�� �����^��ʊ{GJt���ΧAzwU[�]�o��s�#�^���m���$B%�$.�qN�q��e�qv�N���t��u
yt�4��)��6џ�Z����H����9�h��mӇ`@�.���Q�e~:�Ӽ�q'jx�n`�Đ�j6�%ʚ7�n{�s�0E��@�;$�z��,�f�z�=%���=װ�UE/W�6b��)po'X��ޠ�B�'�Ek�sWf$-T��k���<�Y'��[�{��¬Sv!]�����<ʮ�E�	������l׭��w?�^_҆[e��!����u���U
�#�I���G��!xY��X�^/<��F����7��\����:h:���vP��z�b7�=�q�%�A�Lӣ ʸW�����k.�k��8�hN��"10����4����y��[I���9j�2�	3�if�58N��X%X��$v�a5�ARb�:O�u��y���?�P�i{ͨ��п ����z����m3p�Τ�� �b�������q_
fn��, t�Ս��8����x��q[�ƾ���u� }0�Yy��9���	�w�O�?��R3��5~.�x�h���v���'���z��\��\�xg�чRNDG֢� 9]��ri6AD������^z��F��Μ xO2[{اs}���cfUsS�}��S;	5Y��X�+�.���̝b��E������E���%V�h)�̳D��c��EhC�=�f���Bf�R;��a���[��a�s�$B��8=@8Y����v�����+�����oŒI�����>K�7N���W��w��{���R-̻�&�zA[��"�;y9��K<�Ia�`�*X�B��U�c��4�}J?�T��9�2by��5���LT�����Ez�����%&�����L���-����=�r�uN+tÞ���jǁ���-�kwh5\�mC\+]lSԱ8�"	�v�j��>llm��x���G�~n���d�����y��55	[Բ)�9>O��S'�]� �D�xo|r�&0���@��W긹���	p����z�1�!rD{5�?�4V�ϣ�%qXc��������7�L��n��!��"n�:��{��^j�A�����һ�
Y"q)�]�e�K+}�<�}�þ�û�t�
]�R�r�����w�&@�L2B�����5�u�I0O_N��l⾬���~�_�Ө|m*�����xJy��m����1>���#��e��K�������q��[�NZ���Y�|�2 7(�2�F�1�Þ��A��`�����L�+Zg���4�9�Z��3�$ ?2^�L�!ˆ��xl��IE鿒τ��}Q`aBpu����6�(��ɯVL� �#���ύ`����(��"�
Hg��k��4�[��MP��U[���}���3�%_E~�@�����5C�����#/5i���Y<�
� �;M����e �N��֏� 8W۩x���Q��vC4��q����>��@�׼R$�m�O4���Ӹ����֩n������_�q����~.���P1��$n�����xR���>�d�?�]-�+��A��.v#���,���J�_�)���e�qz=�����M��CRD�F����R�k�&�,`��=[۝��{Pp*�&���w�>��p�b��C@��t@��������dR��wU��U"u��=�4���� o�T�<.����2Yx���E���AnӼ<�/O�7&*c���H�S�u)��Τ����a����ߓlt<�V���ƛ!��sD�Tz�ݓ��'����}��y~�?��I۠�fޘ��#�M|l�N�����M�?��m�m?�H���K#xJ0Z�#jNkyM�%��~q�R�|�� <�#Q�� ��G��/Q�J���[a�k�f6�`1��㘲�V�W�,�xO�KZk+&� R�k�eV����\�t��:�����Ё��R	���>E庅Xpw��������%��o냓7Y �k�̹�=~A�)������kS��^W57Vk}��?�����7���Uu�,�}�ug���՞,'�M�TK�R��$�.�KH� *��n�f�� �j���-�E4���������\@���WN���_y�_/��Y��n������ph��4^������LUf���P;U4�y�b��麟�	�Gv����KՆ�0ȼ
#	�@?r"��`(��+���`���gm�m����{���@Rq�m�����-F�ӄ��A��<s|_�.��Ca}��0�<�����-�[��j)�0���Zm�B���|������XĒr���d&"vAA,LŲu�V��͆ď��g@��f�d�|!H��]*u��צ��֞�!���g8x��}�=����`k���&,��SKO2.6���?٨h�hVg�N��Ǝda-����$~�^���9�,;;��D@��ZpU3��}��Q�F�q}����빒�{zZptN�>r���=�YR�}����8��a;�hɝ����j�dU\-��8Qo]花���[K8����[wشN�e����	��ӵV���	��1ȸ
D�@jS��@�� ;C��qyg��fKm�"��OZz����*��\/!�+<��Pc�EH�t��IۥOt�dt�̝7QP���$.l�svŗ�n��������2s�����%}p������i{i����3Ҵ����D�,��x���^Ͱ�,��Ă��"(��P(k�VW������/�W\��*�Z���y�l���v�Xo�S �}��=�f��,�X�t�c/6��)�d���'�O�4���#|V��+��{G�Fy����^��t��ڪ�C���ģ�'Ӽ}W���@{Z��(Bz�y���Mc0T��l9�&+�o��7�Lk������o��o�,�4�F��822z�Y�~F3M�l�F��i����@�)��|��rC �{;a��ƞ����繋��,5JE�?^���Z�Ϭ��=������mԿ�_��~ꩡB^z [䴏u�c����vp}��I�:{�u�I�C��;T��	�5��ߦ&����K�xU/��9	��d�X��-��ώ����=�1�{)`��?�IK��?��W��Ԫ�ݾ|"��Q�md~N�y�,�&�v~B9��x/j��`��Cn��*L$,�.9t�f�9%��ZMvg�W�NۥL����/>nȣ�ػ�d/Ԛ)ۖ��?y͔�bM���?�S-�z�)ik�H�y�\~N�	$���GɻD^T_�~y����9�G����2�H�II]���X UW�Č�p���+녙�-A�ևs�����VLE�.:L���H$�S�Ml8J�G����õ�z�m�d/���HpA_�lmH�vt=IH҇Qs�&�$f�T�u�R�ژI�T�O�i��@����L���;c@4�^-�sp��g�;�̳�A�'��(�ќ��`n�D�|�v��H&j������W���K������k�QS"7�5v�5�sQ�hp��+�]�0�"�$�1�"sgC�8R(^'�YC;y�(o5/?�khbg�U�ŀS>��	0�`,�xj\��LW -
o�gf_�o�������u�q:cq&%Y�rr�qQX�(I��BBb�8�N�y�̴��L$�v[4w('�FMV�?6�e�7n8wAxy.��G��2^h�Qt�
�6��O�k���������_p�&˖r5ㅅ��r[t�Ӯ�zQE%M=���e*�0M�״_V��]а1TѲ�bsd)���A2���7;�
�Fd��P����60����9Ցc�o�ΎRh3��9�{aA�PNa��wy+F%:n�`�b�ԝ���Ȁ���嗆Q�HD:�Hwxs�b��;�~Tܙ�%��r�����ol*O�(�Y�*h����?��CK�Y]f��ʜ
�5�n��q�ڀ�Һ4���� �rz�HO*^�X�ۡ�뷄�e�M1�͆�9�"@{�{�������K{j�@W�|��)i���,r������si��ܯ)�z\{N>������S�_
��~�<�h^�&�4���P{N�G#	�k��	p���d~��{��
�_D#�-��h�9�:|���Z~�\��*��g�5�Z����7�$Nu�+?g�����o�kY��Wh!7i��b�P�������
�b��Y�~���!N�Dx��fb1�� �jM���\�X�Ix�R%~��� �8ltm�~ц�]�qv�G���z55�Z9ELޏ�7�M�Ԇ��~2�޺z��>\��-�Z�Gtތky�K�p)�%�3���]3bd��5�2�-��$j[��W���(�Y����G�O_��L��g�
e�Jص���~*�'��^�D����\�i��I��}Vn��lpȭψ��NCn���f��k�T-j'6�d��*��s�h�#�C�#���k����5�hj��X�� ��V�KMנ�f��e=�4���1��ѣF@����Q�d̊t�gN�J��%i��X�I3�d��+{�Z~��iM�*-��KL�t�N�lE��]C�al|m_�ã�F�X�����r��g�!��$�e���\zKY��$�����ѝ�_��i�U�f�3��������gݛ3�c�7�5�1�5���?9j)�5R��:�lX+g�a�XxI]�����Eۥ�Z�Y&%�r����(R@{�k)�����(0ccRc���SXW����W$a*�-j29~�rZuf5n�^�wwZ�j�m��H�p�d:��B-�5	����{����ҤI�|�±��&�Z�I2 9y啩Dɂ���O[�\x��O�381�r.ƈ���K=�sg��/��6/�+����S`q^N5:Xn���!�_LߕR�M�P+m�����!�r�8�xݷ��޿bs�[8��8(H1rTn!k{IZ�P#qAx'oŒdl���:��4w�w���S�^�P�gC�'T�6SAG4.�kF8��k�=�p���*��X��ɇT����ɨ����y�~D)�mSognΏ!�z�ؠt��ݢ�	�4 c\tB�QS��_l9W��-p]"�I4��4/Y���S���mCK�g#�/����Y|5\D4����i��C�FS&]�^['��!W���T��d.*��X�cl�_C�O��K�q8
�ff��_[
��SD��,����H�,��v�
�"��&fy£�(��*���Jq#���#2T]�=E4+5}��&��t/l >+��vJ惰��n����}��E�z�8�rf�2���wb���_���w�#'l����n��r�2
Rab�� �!��Ka�es�o(��T�tHU��ֽ��b �h�V]W���Y$is8��-S���0�W�V�^���+���};|������;�Ť��[�[$?#�����o?�k�(<����f^��t�V e�YЀb���aX���|��~������J�fQ>x#�N_�9��k�W���rZ�^�-(�)I��0�dx���SD�S�����S���؊��m���0J�?b7� YTx�����F��������_6[��'��p���b`=�#��5��HD�l����gvX�P7[�=M��K8��v��*�(���!Z�����3��2��@�"ե!���SJ�j_�P�3F鋔WY��s����۠���އM�K���s]�}1�I���(?F��"�
|XFW\0LVD��#�V����G��XsGOO��g���ֈ��PDӖ7��KD�P��2˂7�י\4�^��T��!.9��Fp�uD�o-sc��i��PMNz�m��ܶp+m�T��=rk� �b{A>Sț1n�ꖟ��O�ʯ���w��ǐ=ki�-"Z؂\�)�6n�2��ZL����+W�zg�ܜ~^T��0�S��`]a�����C�υP^(��UK-��|�������9o�\��C 9���g={KT\K�#u�˒��'ח�=@j����D����J|�x�>%h��|d�i�(
��|��"��3FmOM��_K�q�׭�����']ݮ�C���隣#y�m��ƶm��ضmml�����f�m;�m�~����9�W����U�VOu�����,��\Vi�������:�dz�P��P�H�/�dr��X=�8�"U���Z��I�g-�e7/�Q�RG<�&�P5ev:>~x�E�n\_�)B�Po�*T���I��H6�<u	�o5o����T�Q![>\�OCu��Z�z����I�耱�j��&���&]D����L�
�6$��t�W<NoMՔ;����bcǭ��GMy�<�MѬ�D���,�E���L���RNLJ�}ɓ�dhb�W�t1/�Ǔ�~C;f�d�M�V{��7�P��е�	"�Vk��0�BJQc<��wV��KA/n�/c��O��Y/&�o-Gfb�K�*�VHE���]ƗN��N�9��$�/B;Z6����7.Z��H2L���"��4FZ=�@��b�����)���&E����/\t���%t�5|E�����Ɏ�s�wʎ��ɨ�
.Ҍ�td�[�,u�Z<�� 2�?u���FJ��lE�MuЪ�,{�8��::��-\��1C�j&Ud�cV��R ��J1%C�P���Z�o�dT��S��tz��n��d���ҙٹ{����[� �w!���<�|�͘����C����krX�TP@�}��Λ�Q���O���wk��-2��������[
7��K܅̵%�y��C��#R��akW7܅I/F���A�b��
yd }��Ӝl��}M�%� ���E���w%ز���y���ӄI_
��#�V�yB�bTηN�\ȿ~�G���� ǥ%���YE1��td��ܽ]0��&�N��p�7��[za�U���a���'W�$����-� .��:���y��~���?7rtǥ�VQk�~嬫ۥ�=�j�ΟN������*��.;dL�ˆ��͇I[��\��-rדx"��=���&�k2oO :iU$z�6�8��r4/����Y)����y��T����8��ݡ�̓J<���/��T��Sk�Ҍ���W/pc�%��>R�Xt��3�	m�N)��^�a��h��i�W�?�n%W�3�154[��6�!�b�L_>���#\��SF:J<�o\��2,|�$e�,z����L��c��v��Hx�cKҚST>�[{s�oF/�T'ÿ]�(}�_�bR�����M�[^�Y�HHdX�x�-������������&�,Ɵ��'���q�����ܺ��J=�?)壮�M8����E�C�P���*��}�l���:�v�bst����#�����N/m!ֳ��!4m��"���b �AO}8�IGc"���̍��tsvP�]l��Q����&��⍢���Q��,tNG��xx[���M�L�͵&"�:T����m�0x�m%�l�=)2Ou���H�%_<,�~��2<��s�h��q�+�G_�x�j��L��>Pf���µ�QB{X��҇���4�b�Ѭ٭����#Q�'HO>PLJ~y\�dCI����p���s�p1����\ge,�go���TA��,"�*j�p�3��/xN�"-&&u��Ů��'tO5V�j�2[h=�l}v�
��Y�Tku�wvX�3x�)�I7�'�wo}�y���/�?�[�h��RQ�7�j�d�8��!}Ƈ�PX���B��9�vvC��2��
0ф����m\���vlκ�q�rX@~��6�qv^�<�+�Z-9'������G�@�A$c�:���H=��-���.���f����6<�esf��i�pW����.������	���ȑ=ˊ�@ ���ʝ���6�X�����&�q�Vz�F9�b�������uyٶJ��u]���&��9^��,O�����㽂�Fnk�s�;}>���s����c�`�!ZL�4�������?� V���|L��#�W�Z���l��̼��yg��1��Z�z�G2�s	�@\@��U�[)���W-D���VT�	Z�����Z���*0Kx����?P�V1q�[)s��>������-2b�ũ�C��u��=)GhqJxkd`2I��wŤ
ma�g���v�md�u�S�֯	�L��?pv��&B�xٚ3��v��J��l���V��.����հr�|\���L���]P�q$��ߓ������o�m�C%�5i(�=L^��d�8���=M\���{t�'��:���{hё_+G��}?�J*��X�Q�o�����4+�\���1����-VMԖ�wO��[�H�#��/���}w���zv�&$d�f;�����bS[b�����&�Dbc���O���m-��I($	�`H�}�:76��q.Z�in��'x=/�}��'_�Ȥ������w��ȁ����#ЦT��J��D+^�8�����o�WT$��(���$�C�j]5M/]�)7�Ҍ��w.F��^��ŬJ�~}?mg�9#��aQ�=���G���a�JS�2�?��*��5AS:X�	i�i�� ��3@�eD�Eaf����!�*�a�����r�\��wS�A�.y5����#F����d�y�bS^�x���@��DMu6���l̞��-����[�v��U�"u�e�O<
W뱼?�-�v��>�K�9B�`��pv#ׁZ�%3 C���J&��i�0%5^�i"c��B��i�d�PD�p���U�L��ou��c�9�P-�ǅ���U�]ENn���O12Bu�L���[�yU�^q�9��#,Nݜ#�{l���@�?��������j�٢;�B�|���;�+��2T�8>[J.F#��
�͟�v'��ÅH�l�AKuWh�D��?������F� G��ld�O��
<�H�^M��I��@<�E�������9�l����L��'Œl���J(s��7���RY�@�<�IK�Y�}������-Yo��QnB�G0���vZ�[I� 邿��b��Y=�e�����P�`�p��I���rd�o�T�>肾<�_�h�$�<buj������W���~��т�6S����ErX<v&�U���C��t�~�<O���_��\���dȞ����!󶱼-�4!�߈�R�hr��t��-����ߊ��RNCz�w3F�1g��iٜ�H�9rҽ#c�V���ج�+����{@o�(lh�=�n�h2�:�g����͓���������[����cmW�C���$?;+ m!25����i�>��-�Tp�Rh�ed�]o��v�Y�P��� &9r�i����5��,�<�:U�R��y�-�g�f�ui��p�mo� _���
F+���<�xO'O	8��)S�
��6����ҕ���c챣;�q*k��V��8;w6a֭� �D��ct�IƄ���(�и&;�a�O� ��!Ldn�N���řX���a�����.�G�&��ܔd��r&�v�c�iav�m���~Ǉ�oͧ�*�]TD	s�"'�N@M2�il�yG�L_#�o=�d�43)g��a ��f����	��U=�b�����=
c I��l�4��`�#�@Сgܮ����IOhF��Oj�3�&�?�fe��S�?���~�Hl���.:��zd�T�h��0ڰ�>��2��Ej��l��<��~�lr\���n�`�I�����!���]�
���,�A��4w	��K#n���7����JU��5Ma�ͻ]��]9�����\w��S�,-�_4�f��M�����:���3Uod�F�U�m������|��u!�y<����Oď��$�b��,X���E��q9��q�'�nO�Ŝ��ok�/��2)+�-�b�u�N������"���}������>"��u*�}Y��z�'��gew��13Ae#�]�@SF!�J��L��͡��X|x�Z!��-�vP�d�)_`�{/��8a�Y��LL\蹑�':2?����	#TAD0���*bI�BY}4��"���`�/�6k5~pv�9g��v�[�q1���K!��}|����T<�{�gOH���Tz���R_��
ݗ'+�����д#��^>�> sn�r��_�R3���0����6"��,����Ë�}R����I����]�-��iH"5|���ˍ����`j뽶��7�M��?���`�7��21G2��8��}� ��sB����c�c9~�UY7�[�_�����b$ɩ�G�ސ��hV���Rk*�2��'�j߱�]f%�j�N�w[v���=�-`�[?��'�!�>���e1C |R�(`�>a3'P�j3o;�d<���]x����K�bo�N��2�ZRB

�=
�K��f{0���'��f_M���Re���vS�O���}y�z�~]ؚ��A����6�Rkw|�f���J�~H���|�����G��\��S�������ʈ&��}�X�w^XB�6�:�S]��bW��S�]�k�us���r8埞��X�'hg�e�ky��^���]�{�E8�^����I�)�cȲ�a'�y�@���n.z�BKٜJ�ʱ���x���ԡl5I��(�t�[��$�U�~}6@�C(<�k�{4e�i�p9�U���k��j������=�[	k�B���v*�#����+�?��&����U2Y�;}�kB��3�
�Q�s�F瑁�&ͼ��T���DT���Bv�!�����ǉQwʈ��O2�A1��	E.u��:9��]���V�X���l��/�k_��w��4��4�J^��N����Mк
��Ce�8e4_U���\��u����X��r:�q���Ӑ�\45�cI]﫳".��:�� ̆���@��L�*�D�eTqvb����Uǂ������e��������X��:vu�}J��S�>�tH��?	��7'5�����
��Tܵa�ڶ9�ϟ�@�R���>��]�q��|wjk�#Zep��147T�ڰ�9�����s�s���(�uܑȒ��̼�cYy�4��J��ΑV ^'$�Σ��Ձv�^����A�������n�������2iz�jd�h�/ ���г�����z�viNϖMf.`��`VWV&�Z:�ovuR,+\ج�Hٓ(8A2�����k�_L0Y+�6O�Lo��Fj)GF�kF(r�_3�k���u�)�j����){l������U�|Q�NQ`���5_g�n��Hj�r�������N*��?˧d�N��h /NƮ3��V��vA���d��O�q�+Z/��{����K��dDvR��3��N�4�ZY���Ѯz ⭙�u�>��˔��z�B�Y���p��__�#>Ө�1e����&"Zi�v����G3���8�p��9�l��T�{��,�zu�+Ҧf�ԮO���aM��Ar�m�e��vJT�p/��f�g�we(��O�?J6f��|ޟ��,۽u��<gJ��I]�{�X��>���j],>T4M_���Ji�c����?������~�����Nʪ��Z�ib��$�Q���o`��V�j
�t��GS&g� ��݄�x:��ב��������O�����s���38���v�{)U����׫��Zò��N
��K����l�?)�������'
0t="��!�����?�೶���	�'�"^��Lm�H�9ʋ�X]�f��'�
��ͨf�x��D�ke��ڈ$(pJF>w���ΒE��"t忾��p%0�׏M*/��3:�]���4!��"+���L6!ʿ��.�L����U̥�Q砆`/|w����hT�u�8z�c�o��JL�$�C��1�p���x�i�f��8-��n�	��o��A;�D�H��OL5t�]���3} �<�Ө��0:f�n��=��)�c��ٔ�Υw�ǃu*פF_��n���OjG�WK��%��l�3Ĉ����O6d¨�3�+���U[ZIy��|�`X���0lںwqu�v��}L	p�8�9��i� _�����������ϫ��byi#�,B���2܁g��\�ț����ݎ7]�}�jM�l8&���vB�|ѷ�'��#)41p��L�%h|���]�s|�KEs$}��8�
&�v+c���\Թ�ݷ}���N
�ٗ��?!Xx�:�����E1������*�>�lf!CSE	v�!]M<�Yy����ӲԆ�>vv M���Bߧ����ٍvp다���Zyj}v랕�7 $��-�#K-�$� k���T��:����g�u"i_�_2�>>���<j�w%n�7���Һ�$qD$���dN�V�=��v.��L�ߪ�5�.��#���D^J�Q�:6���I0�������lܬrӜM���b�PK;�Wڂڂ�ڒ"���9؞y݌�1p�YبO3�tT�������6%[�Y�ޭvL�r�+���h˿��@�Z	�����u�,�!k��d�h�ٕ�T|��`��+t۶*�O�ؠ��^Q_�} ��:þ������yq���$N+�Zw�#�jt.ͺ�av���Dv�G~���ۥq�{�-?$P�/O��u���s�V4�#�Ek�T�dm�0^�ul�!���V��J���Eצ0b�s���(�-�8o��k��_JZ�y�=�k�1�hˬ�᯷ZA(�;���Qd�k�-�K���~?^a�U�S���+,�.a��m�\����-��M��������:LV�7P%J�����C�k�>�9���|�S�j�j�}���<�k��ل0��0n��#{��;I5���nDͧ'fֹZkZh����{��e����w���V�`/�~���+ݬ*�~!3���:Q:!%�UORF~ip� DO�*6�oo}�D;��Y���C�����?�
= ������Ei�t�7:�o��z��"t�1��,�4X� �ծ�v��)#�T�'�ں��ҕ�ũ����Өo��Va��dy7p{F1�u4���4�@m��>~V��}�Y��:��G��"?q:l;�Y5R�5��4���l&������u��k�ʃ�j5,���B�LJ��d;c���!�n����5gAs�6ʠ��(N�op�nE���Ƿ��2�oi��j�Ic���}0Ш�<_�E� ��;��ď���?�}2��DSp*:`g�oh}����Ն�S���d�q�V\���O{#P|Wf��g��H��:��8s W7T��V׆�ͅ�Í����݀�F��s[ 'd\��8��C���*��h�����K���<�{�2��p�#k����y��/+�[�]ܳ�(�m1U��[(�a<f��e�%L�2��|�m�s�SƈE������ ���V�=;��}}g�R�����Ke�Z�߽�D�@ϙ���z�� �uV?��7j�+�.MC۞'�6�t���tR�q�~d��3��EFq��~�R>m�F��*nI𷱴��w�R�֤��������0�"I�^<#��y�>��P�֋�5=��TZ�d����5x��8�V-��T@y��Gu�t��2�����&9[\����A]����LM�]�=�>�ǿw�b�N�)���7�U��֍b�_w�è�FRu�?h�LHҿ��y&q�H���'�Q@;�*������G��GΏ��Lڮ�%�b�a��q���6{��u�b{����qC`�e�*4�$�՞t^�ԝBg�6����xӜ�� �o�� 4�tB͢��d&�+�+
�&cF�E�z���z�����\(*�@ꪀ�Q��u�C��p�$��5�����l��XS�3�V�F�����jK�[ �`�1هϨ�������H�Hh��i������5�% ��ᄣ��,� 9t���О1�g��u�Tm7NaW��esj�Qq�s�����Q������*������'�߄���~����|�� �f}G�tXP��4��*7�S+m�E�,�K��.����bVu�7��itG��D T*���da������x��फ़6V-��Ͳ^��_��2�E��4���oۘ�y�
T���6�����{�b�U�^^|�:��;[�
Q�3'��]�D��`}�v�%��z;�!�y�9Vu�Z'��T��(y�z=�\"��7�o��PZy�[��\�I��z^����0~���,�$��r�5��#�m�qM�U��B�%8Қ��M�����ُ9�@��t��ì?��<������/�.���u7~�C���K�}�����)I�����V��s/G�� ������=�%	����j����a���4���L�g�z�0Lr����� ��J�����A=�v�3�!eSP�zOj����$���Q�����%)��Q��W�P-���?�[����ץ8��Y�G�ƥ�c8��j5᜞��V��\��*�ƂkRQa�s����;�Wo�F[�9�2�(�"���\��&M��Ѯ��y���ӃET��$�6�QI��	���F���f�4��"�j���|"H�x��LH���~��]��dI�-�����oӎ`�MC�(��AF��=�=�
��������ա���xϰE�G�����rBڜ�D��Ͽ�.��l����1�h�Q#]�����c{,��4�̹Ȋ'E7�w���FT\L���n<[�����T�yi���@�q�s�ܾ~��{/.p���bpƺ誌�6Þ�V ��'���]o���
!�[H�O���1�T��C�f�(��4t򤟖�l#�+����wtX?�K�b'���TqC��[���+��q�׊u&����HX���Geʩ���ʏ�'�y�ж�y=y?0cB4�=�@ԅ��w&t��"Z.���M�
�+_!=�s���&���h�VC����:�h�a紕����{�����0���� mdB����D����5u�N.ӫ�)E��/n.��	S;��Q����XI!��.`�
�w�Ç�l��7 ʫu^����TdƎB��0{PoV����W�[�3�1IO>�ȝ�wZ/�
�����l2�ȧfYK�Dz��kƻ�� ���DEp6�:oZL����.Ls��Fy#��̘�k$�m��q�뭮�:��A���Z&ѽ� ���9�J!j�@�*L~�e*���A�1�L:pk�����?��Ʌ�hϫ�{W𾏨D_'���sPr�n�f�3h�%��x^��۝�<���Wc���Ζj!���1����>~�}�/�v ���iL?��^��G��UVxa%H�yu�:~����qZ�m�6QSF�j�~��o `BWQM�Y�Ļ��~��&�����@~��=�`��	��]��|�*�|.[-�߭�5�qf���颿I2��pM�	�s��
��k��={5A�"�T��aq3�o}�ka�w�B�SM��yt��u��I�y:�d��n�;,D�Ԅ�V�?�����?���:reݟ.����(��$J��c�v�ӈ�-��q��g�Q�sG+�`������/Ɔ<#^w-�9hs�D��|��E��x��'�ǭ��ͪ�A��;ҧ���63����kwc2��^�1u,Zg�v!�J���*w��%��cƘ	��<�"���~{ʵ+����Lz�lm&5��w���EK�_茼�{L/wM� h�;�-�ŴoW��	��zP���ڀ���O�
��M�^9K_v=:�Ƃ����f�~_Cr}P��ΗSZY9RG��ZF&�����LL��ml�����!�3��YE1�fV�G��!4Gyu�/��Q�%Ly��-k�V�YO��ݴ��aD�ClDR�rs��-�G_�I㶦��/�&^wex@�X}��.Ea��lC:c��&�`���5�`j{V���F�M��kI�ʾ$�D�d_����?ZGG&$e-���X��¶���+q�j��]�n(vf<�v�
X/�@�TE�K�g@_��]������Z�����9���Z}� 5�u�u1Jq�'�B������X����+��B�<yrt���>��u{�j��G{|Pv#�;<(o��ٗ{�f������8����ݷ���U������(�-	�a�<�.�����3�<ބI�Q�: 6J���}��O�"�y�g��u����lۿ��[V�N�F����=�`!�O���gqՄ�����@
`?�7ihj�?܃-~g��(��Q=�����B� 1���2��=�aV:M���������E��&�k���G�W��P��܍�?J��_[�X=bC����H`4{�0�0���\�p�H�D�>Qc�}R@D��+�`8�`Z?,)v�?���C�8nU`��q�!���@I!I;�HM�*?bE^Hs��5H�E��*/Ϻ�&���v樎lmC�KFI�;��@��y+������Ї#
	fM���F�tϢ�zNdvk]P��	��q�|fI��W�:��Y2Ⓑ9@�E;b�gH��dA�c�-ޏ��2�����K�Y�!�S�*YM�ЦU>��͕��"�Ou�k�?e#���i�f���Z9��J���0v�)
���UB���C:�ѣ�^��{{��}�^��>���>�g��Bj{��yPR�@��dv��{K�)�A���ЙlG��Q�Ƽ�ss��q�蔪�e��|�J�G�Y`f0�20p2�\�pLXgܘ��Ea���f���^�P`��My"� ��C�K92E�D���>na	"�~9����V\�%��c��m0�&���Ј?U_�֔,� �481z*So^"n?Цl��PI��8aU��`�k�}�+4��ت��`��!�Ĝ>X�7���l���T���]}�EU���ld�1�Ty9g�r�Sjgn-!�);�Q�ԩW�W��C�q
�&s��%�_�����:��9���Pa�O��$I*O�hn.��[?rڽ8�ྱ��&�zi�����D�r�ֆ,AK�Cc 7���j#��9�RPxo+�,���r/�쪨ë�YU@���Jp�`��|$��z��A��3���٪��D�'勘*U�����D��wb��k��ÿ��J��,��)�9}��rJ�/�"�E�~�\x��+m�ػou=-8��F&|I��*!���j�(���#Ī ��*9r�sv	�1Y��c=�P����LU�Gd6�1xYrLZŝ��5ءd[>�WhV���Fi���.��'&�TRA��C��0�5Fa�~(���b Q�fF�6p�(�#���#���rb�U��qް��DSΎ��9�7^{�y��dˢ/�s;���c���vݤ�J�¤}I�Co��qF��ߦq��v椑K)&nq�]iM�T��+h��?�}(d{�U�(����A
*��Q/M~Ņ��Wn�]�f��/2O%�"�=G��a{M�;�"�U~���J
�?ѳ`a����Mج_xPh�T�2�~8ﺴ^�#��8�����տ�H���J�/⅀_��AJM^�h�^���	�,&��d�j��:#�D����T�,�n������r�ݓ�f���;ǉ	�.ܙGU��?��/�ɮ΁Gj�.��͉� �z-��͉�D���@/�-����M�sz�B�g�+��������.a=����;`fY�zoM���M?�}�
�/��T	k�`O����sNT1ic��gC�G⍋h�5:�ٷ����+�?+7=��P��]@艐ZA����O6�Ki޼'�N%�V%U>_��l�E��;ٜ�I�]3yJ�r��Pt��!����_$+��wC�{#�9�8L���p�=���Gq?�P$����ف'Vv�{�%�t�>�à��*bzE��������j�3+�����&�U6~_�����h��lw+��b�������B��H|�'4�=�����r�9T��Ʀw�����ys紺[�ۛ���t�q˅]l0�eiC����]������f��~��3ǯ)���e��u	8�����;������O�(��o-�\n,y=��}'H�ļ�nI��i��8�E2�af�
Qs�`�am	��cn�)=ۇX�T(��Ԛ�@�vI%�/x�t
$�(���^A��Z��͉�+���tgrLx�	�??���5���~��:;QP%�$�r����~��K}�ϛF
�O��"���R�-�H�,3��|��ӆ\A�����Z=��/56�o�4Q�uw_�Um�d\�L�-����k!-�?v�6�5���]Yw	P�q�&���Q/"c1Uh�;oAxU�d����d���{���+,���Jn��SFǼ+ښ�y�c�6�ٞ\����_T.�l�HS̆�p ��ȄX��#��֒��w.����~�d�j��3Uv �ž�G�&�H�r2w����+����2��$�lژ�:a5��'~�;K<!�����Pk>Nj�jzU�W
k����A 4�v?2�堐���=��������9��6b���@GH	,����� ��SSp��PĿ���`��V��/`D3�b�����]�a�oUe�	�lc���'�K��Ζ^6>��K��F~/��#�y�jm������r
��CA�|>���g����fJ�
P���8��E����
�l{�#Q4?"��%{�Jבd_�����B��ia��%�9���Ϊ!�Ɣy$�]�e�ٖ��K6�.m�������zL�y�cÎ��a2�����pl�p�~u��(��ټt=J��',����-�=I��{����l�B/��P��5ޚ��g���<�^�%,=��>Pp%v�d�v��:�]l?�K�F�ʜ�k�Y#NdX0A�{�J����U�ZL2Akj7�dl�w�Ja��ق�q6>����r�_Oϱ�Sy����8�,��9����T������u�^:�/ ����wB���F��*F�xAP�'�Bq��-��Td��_7�����@���dR��+b��[8f�5hܲ�'�� w²�c��d�l8���ayĽ.��m,�~Ҽ�v�W���&.���b�W� zypC�kU�3��N<���/��e\D�T���.��r���B��Gh������4���C���s���E���à-��	�
Eb��'��Rd/*>��`�a���o��1.M�'�Q*�I%����Y�Q��=m}�n@9)W�%�N:pލb���w�I��׺fa3+Q	�xHi�-zX�Ϛ�dr�O��C�Uڜ�$焍gn��N��l����&aŌzs�Ŧ:�s��"�!��ӭ�R����=ܴ�.�N׻��m )���k9�8��p�b8_X|�Vy�W��A\�q��;��iW����
i'���b�<Ԓ�Z-ݿ��bc��ECU��(��5*�|�ӝ����u�+Yr���
������̕Dð8mmr__�#���'�/8\��� Z���nN��)�>�'f@�݈i~'���@�JA#��P�_PI��)�'px���b�h̪
8���^Z2g
*���ҹN������e��ơ#�K��]#�3��,�I��r���n�(�+��͍A 4�m�VƦ�0%q�a���@v�[��h�LQ�n�Z����M�
n`]�W&J0k�2c�#\ۚ������_�Lz���d���e��H_�d�94�?�=䩒w���������_�vP��,ਔrc  2�XI�/V�ZQ�d5�K݁����]/FO�Ջ�e5����7�؏ƷD�@��/f��wp������v��}+�P�!�V��~�����/���l˳��
�X*�¿H��Vw};;�?[���m���%��q��x���ł5�OKs�2�Ц~M5�.Ч�ޞ��-��ɣ#�z�����;��# ���{�(@	̀n�Z�a�ZqKx��:�R�3��7��H�Y1�%
�*�y|9KL�ΰ�Q<ɘ�A��N;�ݜF-�,�X2�m۝����̠N�ާ0ˡ��5�~D��5ɤ@���ɯ��b2���:r%F�_������Ȣ�?6t�L��:F���E
k���m^+^��;J�Q	?�yq���?v�;�S`��C=E�FU���!�X)��<�:�!�e��3.l)�:t�92j��0�灏9��o@� G"]�K]a`V�_�a��"��V�Wfdvm�, �`V��E�`�:��'�4�����Z�J�t�������Ӹȭ� w%��*zx���#��jpw���>�[�Q�5�.��.�1�+c"��U��s���$�<ʤ]ηf�����q�V$���(δ(�`$-u��9]ID���B��;8��Y�7?M
n|����1�p���g�����c��� �$K��Cls`�x���P"����������D��Z�aȧ����>�K�>���@����R���Q|dt��z;�|'J3���z��M����lٙ\E��}��$+P]e�z�,6��b���'�~�(�^،$;יU}zaQ��_Zf6{��ۻ[y�U��0��Ef��eoi� ��_��� A'�ʂ#��#t gl���DkVW�/=,`��w�#Y��^j��'�e�a��W�TVq?7�Y�v��2�ر ��F�� ����b�[,���?�⾱��r;}(��7-�F�Ѫ�d�?� ����>*ab��q;�u��Kz�+爗7��T�UDk/��p%��U��,=a��5/׏��rǎX71QJ�&9{�p��̻��#�)>qs|��l*h�:�oLcl;���m�1ciSzX�.h{���N FJAC��vx?��D��� ��V��	��&�K��wƊ?-�B��+��7~����x@���>�F�ɖ$t	"�I;��
]/�mZ$"�<�T��j@G��2f�B��D��n��2x���wlS��vTec,�3`-/���j69�	<�����"-�I���̱��t2:�k\)��(���K��͒:���1����~�n7�T�Y�L�`�,j�/ÈC~��j�Mݬ���=2�B#~g�����K��L7�ok�1������@�\������f��lb��I�.�L)5�᧹�v9���J��z�M6��H���N���dr(0����αΙZ�ɿ1��Ə���u��"&�~��bZM;�&�]�m�di�Ao���N��,U؏gif3����͈���{!!�Ȑ��|9��Pa�#�G�?�j�j T?��Kv�>Χ���EIP���rrb>??�LN�k��������)
����)O���b�� ,��>�%���!�:�Uݖۡ"�.����.��D�vww���"�ga��17�iG|�4��-P��[��M��mNF(�:�p�.����,䄱M�m��������Ε�aT��t�4�~5�)��dc;
�2��O����0ܴ�Ͽ��p�Obt�%���A!�ƨ�I��������&�AŰΉ��I��0�`�9)�E��s�>��V{�W���\6��g�>��#ۓ��{���*���,��M��1��dB&��Jz��Y-�U��f��	L�#.�9��C���Ԁ����%ċQp
U%0e(I�Ɛ���1��8Z��JX��{������'͚�l�?�����p��K��L�,�6[ռ|m�".����,%�s��;c̈շ�4b'��gM�#�(�e��GP�y�HO��ӏ�`K��<d�4tU�d�����y�Y@���~֞����[X��H�$@N����>mEz�R��G�e��3�M��F���(�l��,���!��'���J��, Xr�)%�W������5��lD��Q�����u�K�Õ�L�]�v.���H���f`JtF(2�Ӈ�G� �>�h��﷨i��}�u隷1�'1Iv���ks#��l�uÆ�^n���ǲ7��NTv:!ž�E���C�H���ְ�R���/:]�C��oLSx�0�e�6�����2]W$}?ibŶ0�G� ����R�*_2��L������4��eqۛ�EX�S2��vU'G���WyO7ۢ,�Hދ���gO�(��<p�70�3���H$T�a��Q�!���c��rJRӷn%;�mk�G˜/�04����J�B�m�6shɋO��=>�f|0�3ۏrM�7�l�"v�S�b�vg�%��bo�3q�E���Z�F�8���պ��?o�!m�Ha��T��� ���v%�T�3���	6�Q�:rJ5�0�.�v�zSPgju�;�ݎ��G���U	���J�b���Q^��F�Q�-7̬)Dd�̼J������9� k��������rO��m�
���V<c��l`y��%�ݷ�O���8�Kٞ���`�`U��uKyufM�5�D&)��hm�b����8�UR|T���*���q���8Ɛ`���?�hUQ����.KF�a�����aы=k%@�̀�LX������m��G�g��8K!R8�yw���� y�Wh0��ݏӮ���KiയK���8u��z�=-��=B_����&�53��8��K��4\KQZ��2�='��8��Om�����y3��� }����\�č��MogL<T:_y�ݢ�W!�l�ޔ��w�},M���!^����0�aq[ �[p���	������݂����������������骮S�r�f~N�c���)�p̺x����
�rq�R͂��G�����.�˷���z�n�y����6x����4�~9�6#�0[M.�y6%����z�ʃɕWWM��FE���Y��:��8�T�K�3j'��-x\<��bD��bP�����P6��F�HA����}�A��mҳ{����x�����!���[���ƕ��1r��}!��њa�-��7pE$|\�G*�(x|���ܮ܄/���mυ��`�E�ڌ��-Vt�m���fe1�*g�`߾�W;Uh�gpq�!�B�i��v��'/��Lg?8W��B�s�8$x(�|uK9h��{��f�Nʏ���`9����#�:��D'�[�L9N�mi�G����"$Hj��䈀����ƭ��p�L�UfEe�fB����;�Ԉ��[7����ƿ�y�˗o(�9��K�ޞ�JA��3Y�����B;������s^��������t%gNL����9��3�!�a|A��j���!o:�4���#j�u��_�f�<2��>��-�uʲ���$q���.+
R����7��4�8�z�v�=_H�i?����8�Q�4�6<p��YUz��M�rƲ!ȠA�m�5E�#MEL9�+��Fy�^iM��U�kIO����
a�i:�[%CS�`�e�2�=��J�%֑�W���or��Ͳ�t̻�� ��ǡG!{���*��)0�4�[H�-���L�V��(q)-�-�?Q��ƻk�v{��c���ʦv�p�熼��������	1�Tf�d�[���݌�w�_�ٶ��XM��L^�c���N'Y����\8� :�S~�Aʕ�8����Q�n���h��W��\hV�u.v�Dt%�r/�m����SN��Q{�Q�H����٨5����rM���k�w9��\�w˟]4R������Aܮ:���"�>���4��7ȍ�;��� �= d9�����)2jǒ�y>������/��Q�l@º�_��E��Y>��	�(��G�3�L{ܯǬ��ڰ�ҥ���r%���mH���q}8Y�1>=ďs���a��6�̘�
��BJ�3�+�'ˏdU�$�!U�]#� )�t��.5F��p�J�=uE&�&�Q���=�]j�fT���yl��ti9� %�o.bQ�S�Huip"~A�PtY�>%��a�|�w.��&�m���=ʖ@/�nYP~YPI���!�-����+h�h���[�Uf�Ѭ\��"l�:��C��w"Irx��������94oA�����C�c�����������\M^��������������;p����!5��G��u�!&���y����:��Sn95��K)�]&g�1��������"	�o�X��mx�ߟ�)��>�=�m�6�.6���'ڋ�������By�qU�IZ����W�
gLH���;C�y2�|�I��>� ��?r�10�/��Lͳ*
<A��4ZV�PL��)6
 %���<���j��憧p-�������UpÂ���E.��0ds2��h�߃�����GU:4�-�x�~�i��_��T�&��QF�!ޣD�Y�\���n�����.������(��K�)BL*�3��'�a�f���ʗ]Pm�]��mbS���顿(��������?ϲ�.���M.م�����$��xA�M���Q
y��Ȑo&f������_�c(��-r��0"��U���[��(4�e}��U�Չ���]=CN�/� nm������[��>b�^����Lt7u��XIvCG�<�Ͻ��� �U��<T�1�#orBɱ�d�h�2
(Z[:�u�8m��V0�!{_ًo�C�mC�VԦQH��������EF|���@��hx2tѧ���l� s]y����YЏ|7�FC�=��r�}; �3���
s�|�ۓ>���R@���iS0˥�NE�qi�3jq}[v;��7��_����F���*�*n	y�\3�����l��=�C�~�z�Π�'h��\Q��O�rh����������+��kpƐ�Ggt2��,S���L��Lc�Zfr�=�'?W'�U�o���o6߶g�����cQ6p��H˾�G[��N�UF-����N�|Qӟ"O��H�(a�TC�=A�T��U���3|9���YAyd#
�E�b���W���E�@� ���.�=�Y5�z��%g�G���3D�KY5[�U5/ �1{`C���QrO�����։c�,J���oL��aG��c�"ǆH��/��gό����Q��.o/�*Uz�}� 1dT����<���ϩ�w]}��y��T6.,����_%��1`as��q������>BY{��#��\y���$������;6���{;��[Uڀ�B=}O|��K��^�B#]"|@�����l�����e�P������Ɂ����P��D����y���Ѹ��+���|�ٚ��� ��V{Rj�Ak�3�-�Zqo!�]��U�A���N4��(�F�î�G�~1��꺆�Ya)KǷ���3�#���Ue$xi(&"�Ra�!;L{��h9c���+l|�)�ɈQ�9��,3{�g"�o���Ϊ4^{����"���߳��vԸ�Z�:�~	�Ip��9]�E���0�[������ZT�t�a�?���ا/��\���0���
�y�����Z% ��c�0�xܬ�m�R��{B���X�vK���l����By��v���(Fe? `�Rw��r��CіP�$�2��ik�zC�{P�)f��JO�nMm��\��⍜E����sdw%�Ѳo\���&
�KEmC3|��E]�r�dʣ��d l�%��a��������w��Z�G���?��\ω����!r*��_Vԑ����>�������m7<�1.�0cm@����5��cq�$�j���rsn��H�L<�θl*�p��x��ɽ�߇�ٗ%|*����R�I7t\�z�)���&%����N���$��ְc�g�E�!Uֲ���]�G�b���js����<�F{�cN ڏ�2��O \|��/�Z�w�r�pck�%���
���l7��r9��%uɘ��-U�ŧ���6.5�hD��k�P-���_v����4g_"�@&}[ 5T}{Ƅ)txXl��!00p���P��7����p�f�F5��:g^�G���߻$w�\��o���D��5���Ĺ��ʶ[�Dm�{�,	ǬyQ�Uޑ�9qG�=mT~%�?5����H�O.��|���������ׂ ��[�
��B�4�;I�e���J�}af�T�ﰑ`�:�o�lO�j����'w�M@����sL+��Qp�.l|����7�u�s�R
�ح7��M9�?溯��F2�BL�
E�G2�D��<�������mW�;�aU@f��a��\ܭ�1�6��ޯ w��ţ���$��$��x�cC������FZ�<�9�w>�w�L=t����:��\0gח��@ y�5��1ː�0a|�y��v$����#����Gx��1q~����{�S�J7Z�(�EH{?�Db!�sm��:x���{.�qu�������J~Uu���Un�=k�������ZP��QH�����8�1NL�md}���-����cP�D/�{�0����	�|���o�9"������E��n��h�֌�Q��3[}ܹ�w�`��g��j�l AB�0Ӻ,kLVd��	f��C�mw��Z[��0�@�r�!��w� e�x�5ʐ���S\�DI{�C���:\��%� d���S.y/�&�~��L*�~��0EUwYK�@J��s�W��:(�⢪3�T��u��cӚ�j�ӕ����� ��+�"	����[z,�M��Y�ک���B��mê萫��/�ɓl5�&�N]X�߅g��� n��r�آ5�mw�bK7 �&�m�|6����/�v��l!�bR��-��0���e�&�`/U�~��>���2�gFc6ac�q�ir��pg�x; 8���,Cm��aP�9W�h?����
Ю�?C��ϓr[���l�T�0hskzh���E�����L�(� j��ve�S�����dQ<q�&I�~	�G'LK`PQm`R���u�SǲD�g~�Q�x�[��0Z؉�q1LM�E����/19~n��g|,k`׸����q����A�
�m��݄�|��p���h��<&�_���#����������%�:o^M�}>��'��"�9�so�zf�M�3z?�SQA�ߑ�Y�A��]�=_w'��P��S5��B7��OS����/����/��$s@���}�����М�/3'��Ȍ�ǁ:c|��=���*�����?s�V��zc�lQj�)�0��ߞ��J�_�JB�X s��/�g.�낐����	�햋��4��~����DpY�-��9a���^��F�
|F3��,wq��\c��N�T��7<?�IZ�i@c��&���s��H�A��^y�VZ�5i>��$gP����3�4ppex7t�
dּ���N����̌y�i.�o�/;K��&^�QL~
�]�M��ԅ�W�Ge�X��F�*�uGlr�f`~jԹ�=�:�ܫ�I��̡��!���o	�n�VEAU5� .'�%WZzPPW#S=J�gy�4]���܆����O�I��~kT8�(J��̮��R��a*�:vA��{��;};{b�E��-��{����ޯ����y��4����n��ڢӄ�G��(���Ȝ=L�i՗{1^Ј�(�D��_��I>�gmݮ�jU��m��3�g���6鮙�؇�,ئ	VRg&�&�8R��mMːz铂��-LG��s�.���wq����j�vB[smq|�����S>CV� X�j�58&?�:J���o��Z�;wޑ� �p��������LU�,V?���k�	��B��m��gI�B�Ǚ��c��0.~����L�i�[MAM-�����Z�=�Q�S^��Dڟ漣ǆ��� �@@o�A�<ܙJ��_	$���x��م��Án����,zM���xgG�W�_���R�@Fz6H���	�����V��X�/(.�9��R��������h.�P����= ����2e��<:{��5(!�Ņ��e<V}?�tl�3�u�>�7
���l\\\��;,YK�D-��~������`���a��;�?b����l�=8�Z�~tBr]�ߟ,(8Ԣx˕%ܣؐ`�,A�	3=23z:�ǳ�}f���_�d�Lx��}���k�H��|�Z����~���� �����Q�I�JoĆH���F*�x�K��l'	�TvXP���c$��;k\���9@*N�n!c��c��D�6-���U v�(N�W���\���Ȩf�W)����ـ��n�2c���Jl�"z��
��u30u��$�ߞk
����X:ձ����Gj2-���S�QSA��UQ��h��ǫڈ�{����I#�|���$��H�01Km��t��F�a��.G�+�e���D����!zp{aq� Ҋ����*"�E��h/l(tm���:�T���scY-��|V�<?�.V��[N�fQ���'�.a��\�4�ǭX���R��^�ٟ��0N
��'���S��g�����Nl���1�a�$�
�psm;��v��|�\�I�MV =�M���j����N�u��a����F[̈3�4(�"�Q����c��DIo[�f^^�c��L���@؝<��p���i�����Wg�b���]���H�q/�C��k�ԍ��,���Y UM�鉌�"�3m2�г���/�����[�Z�M�1�T��4c���TT\w�����~o*9�)BF�0��97��2?����d7"$22Q1	�{��	Ʉ;B-����Sw)�ƿ���@<��1�G�$�;1ⷯF��ȫ���$Pl+�ىc	�(YE9 �!�V�y	�����(�s8D�˺�c������(��/����ם��P��G����%3#0����4hG�Q�f�v��<5"F��%���� ��ӷ7#w6i���#u��‴��PkB!��V�,o���v�L��M\�������A5x؝���Z"a
I��RbDH����B8 �a(S��θ?�9�]9M��V�F��#�8�ʻ@C��y�kP��/�h$����'S=�,��Ix��kG?��P��<.�rA�e���r<t�J��uC�uE�_r���@Na��t�Ѥt�G�y%n��Y���J�	�T��W&\q��r	)���&o�d��V1C�A̺���sqr����{���_r`Wk�`R����
��j���1W��U�K�O���0i�i>�K�\Ɩ:"UX�i+���-8������E�.�ٛ��zj�Zw�������j��ӧgL�wF���Wj�$�l�G���C�Y
_�UC>vj�R+�<�U3�"D��;�`���L��:pxa�A+$^D�3w��_퓟qw2��� �]w�;	D'��T
]��Qr:Ÿ=^S,�^\�B��2�����X0��t��v�cu�Ԯ2w}Ϡ�`���Ɍ2��z���I5��r�x-బj��l+,RrSF�+r��"��b�vZA/��p��+BQ����,�/��PfKN�[+̩�����M3L�#\������
�X%G]�J����¿$�����R�.��O����r*8���R�٣����5f+����ϊ:g[��K�(#�3'j�_I�3�����0_��l8�����9��1�cg�6.��P~̜�Y��g^���A������OA��NUf}
o0W���� =WqH������
�?"���ק��Cf�c(���]gm���7f��g[����E�ϗ����J��Ǵ�"KH��
�?p���C�_RT���k�ь��_X-�{2��WQPPV<$�=@��+�Ë%���m^8��֧<�	�
y�ֱ�9		�vC��ڈ�ӽ�����W�Y���2nڰ���ܖ�N���+�����Hs�Kq���]�gSq�}9�����/�g����ޠ�d�LOOJ>�1��}m����Lj�E���T��oF���M��ث�PT���撹������{�91-�b������щ���-?�'[�aE8���sB���z����U�zU��V"���B�~�_ܪ��i��rU��I���l�����r���.ם��2p�����<�5Mu+e&�o�%JNȉ��>1>N�ə������_QT2'&)	�Egz XƸ!�n}����m�>�,�t�`�7�,ż-X�ɦm1��̾���) У�s@�zN��l�8�������O�Z�t�P�`�0�z���읺��/�'��`� %��\5�X�b�?
[���F��Ұ`@�Y�^��.����1J�mS�����YͣN,�,g���p��UQU�}x�n�Z��'z+�(?��'8��o7cfj2h�#�L��4W�N|�s��γ}/t��ө��sq`ty9(疢Q�!�/��(��Fn���<g����J{��m]-�O���W>��C�\�D_n�;T��s��H�߱=[�×�ě��j,���8s^�\�vbgD/����)�U�n�ߪ^���p���� �ua)b�*+�2��G���2a������[Ybm
'��J�C�s�y��k"ti��X̜�ڨ��\�	�HP�g�14�����w�E{Q��:�S��t�#|?��%'.�|�$��L�-��%����8�G�IYW2�r�F��aTp�X�g�.4��BP�S�w�Z�|8}X	��%I����G&�|������q��hQ�-X٠�a��'�q�iscAD.&��tE��-���c�G:R�v�	+�Mڮ&��32��]C��5b~?�Сy���y���
o&{�S�F_g��)J$��}��t�Mu/�9�qb��pw�q��A#���.��b%��+&{������5�K������{r�^�8i�N�6R�w_�����������=�C���S��P����%��o]���8^ڷ:{S\�n��?���z�?"Y�.9���bۥ��:�/72	��}+�G���RpW�.�@��n�3����ˈ���ǿ��lo�ã��h����ș�0R�H����Rh(<�薞������3����t�i1���3�w���O���%��-�����H�Y�?�-h<��^�9hn(�$ةR	p�K돲��סWy(�S�C��*p.ӻ���ӓ4�OR���������p�z;J>.�^H�+לƼ���l�]����L]-�n��h���ih���r�C��#V(�­�jY|l�����v��L��v��{�;O�X0"����x�R�lU���>ډ=�B���]4�(ɽ���ֺ�a�U-��n�͙\�ܴ����ptW�K\�]NZY�6b���cc�ζ.���3qfV6��D{�z��3m:�Jfj���G|܎�1S^DZ�M����FzyxIi�������\�x���`F�6����$��F��y��+%Ơ��]�d�U��,璖B0��PJ�ա"�AVP~�؅���a�PK��t�i��xI�Uo�XQ����SJ�jMK��[Y:���U��?}���n8�:���FG*�q������ �r���^=��v�c�;�L)2����gh�#3"�}�;�6\����p+��K���11�zW�7�'J�I�DuP2�X��-���̬�V�����uk��z�"�q:P��;�����t�I7f�0"�V1�<��8,���r&���4��� ��n��g�f����<)j�R�Z������HCX�=�*���c�<�9����Rn�aw��'���Jvu�b-�~��0�6�>�-��u�a�����>�������.i�u���w0%���5�/D4xqMB��2�	P$U{Y3cp�!g��/�*^���v�S=آmx���q�
�V1[���{�e��ʁѴ��1�M���|a�\U�U��唖�a�s�Nn���x��{M�yli��fs̛��q|?�|.<\��7å�Y��v���=�9Q��9�Eע̋��`��u���ɲ~�̺L��f��z�_���;�q��0gg�Ty"CAl],T>&K��ő�S-�*�9���R���语������}@|i�h�1��1k36r-l�w���^^�ě�l�~�����B�jΉ�^��A�j<
R��MDt��xL_ޞ��!�if�O�U��v�M�e���U�w�t�U���=P�+��/7v}E�홶yY�=��s�M��gCY�kq�
�"ֺ��D�/��ļ�7����pf�ϻn����Z$Ο(�9?��"쫓�:R�� @k��ɇ��|#>^ьR�jf�����}S:/՛B�9@�:wu4S�1l��S]���W3ӟ�+�������t`�K���wo�&��"�+2`sX�X|HV(S�W�Z|e�^���H���6pO��z94�%9��2��v�n��VogE���l�;��;�(��Vo��Ye�[ة� :��Ӥ]��O`|Z�b����Zfqg@�>Vy��yc	[G�A��Ny�὿.+Y�[�.���xl ���{�8Q��ΖS�~r�� �v�o#G$���)1"h�����F+~q-�����x�;���xpfn�n2b�-Y�
�`�H��0���5��
���- y��.9Hz4�/�)S��l�%���wXic8��J�/��}��K��(c���pck�q��'4A4V"ʀ���w%V�P$/�� �'�?�Y\��x�KZ��Td���]��!����?��D�q�n���X�@�"%���W����@��I\�mĤ���wR3,_�����V��qݒ��=�̬�4���Β��{���/���bWt"H�}���Xs"�٣�6�T\��J� +a�i�I#� 3A4H�o�CL�P$4ᔶ>�Y]Ú��Vċ������pW�}��%��:�<ڙB�%��*�]Lp�|SR�tRb����m]�5Vf��,��� Q]e��ycԋ�����.�S1��S���;�C�&�J���>�p�����:-\�F�����,�mTKu��q�"@��o+���������\���8��W���M�f]Q���8+^=��U���>�q's���ۥ��G7�P�^�i��"E���F;X7Br�K�T%^�D9����.�f�In&�4�\��촴q=<Y��w���MFC��UΑ&J亅�[�XG�v��?-�zu5�H*�]�W�3�ɸdg.�����|�h
l�U��d����=��rܜy+�Մ�^el�J{.r�@��!L��,�D��T;;V��t��ķ����[�/�mE��ߺt�����B�a~ƀe \t���b�b���.�O͹�A�÷lj:��=P��E֠j,ˊ��8������J�Q����;�W �<�O�1R�F:{�F[gaNQ��R��L����&z��K�JP��S������)M\���	36;1��*L*=�>�:��%��
:QV0x�'���a���Z��S)�U�WM﫹y��D�[�b��3NĹ���ϊ��*�<��Z�Xo7&�P���x�"�~s�Y�;� h�AG�
�k ��!�`J�&������)%��}�O�w��w��[;Fy=�.���)��{�r����B�_�l[�̵!��+F�1O�=F��F
nMf.LL�p�]�}[�ܵw�7�h���2d۶���m2;��kv �q0SQ����QK�k���Rb�om��v��;�zZ�Aj����SN(�ސ�\�����^6uX�!�"��X۷��R/O.�ֺ#O��k���ڌ4d��5�%� �@�9I�ݧW���(|�Q��`Μ����쉊G̯�\,��PKf Y�\��^��|;>}]���7���?x,��o�/�K���Qc`"c�PU1:u���ͣ-7�Ĩ$sq�=A���ң{���&$e��)�A��XKbnH�OyE��> ��VU�c:kw����Z<�2��P�8w�a���o.��������Fb��[3���FWtt����N�6r�t�x�s��(totlL�Xl!Hv݅�����vm����f�H:$��wI�mD�C�[�A���?6��n-�A)xH�u+��G�!��P��i'��P��U֗��F&&DY\L��o�'�o��(�k|&MS��_U�q�kiP��Þ�):��m��8k%w�8�?݋�[U^�� ��I=ۡ���xp��\����x0���r�M��և}-8��9Ϥ]4 	�Ú��S~D<�.�ڿ6c���jD���D4~�ֵ�-%)<�ګ��IL�ɧ�
C�J��}�7~� ������ͺ����<�S���U+���#�ֆ����HX��u��F�$u�oIq�'�S����h�<��0�xE�ri	p�+W�2[�0>2��-d��R�<��Ԅ��� �=)
~`%��|Dc��<ɋ#�<��G@�f��K�3���&����bD���<��@ӽ�<�x����������"MX��#�F��$�nq�� ʗ��%��`u�73�^I��ۺ!��=�O��ֵ,<�洹ZC�A����y��Y������js��n�;��鄔� �������k��	0!����;!#��E����$�b�C���̓��t���٪��ّ-��b ^��%Z�@��[�~OB����]�D1���_Wa˴��"5Ș�c)7D	�	A<.Ϳ95d� -��Z�y=��hm����l��p=�'0�8��Ok �QJn9m�_�a�|�dh���\Ń�ܑ�SdX��\����c6� ���֤`9V�0�GM��C����UOO�A>2���O�7Gg�3�kDּz�{���ca̧��3Uro�R��`̛�vLM.P�9	���7�?=�n����( �h;��
^�@ �ƣ�)}�R<�PBz��A`���ˊP��'���	����#wθ��Б����c�p7��r��ʄ�l~b��A+l�4`�4Hu�2��у�����頔_]-�6�{��>օ��R���%=�qm���b7��;e	�?����y[ ���}Z�<�֥�&�v�tno�;7T^������f)/7k|z���կ���|�X��叙�����$d"KM~y-ڹ��G($���/��?i�
�����n&Z m 5(�$8�m��~�]�zP1&���<_�8��op�	u��-;���3p	�P#)m�P}n��أ������,i�x#^z?�6d���W��t��`��O>�Ky��^�F�h�B?;����*�
W_�v�E����1;�S����o��~�++kB=����a��L���!�٠��lD����?yKV��U�x�ոX��P@K������|Y!*��g��!/���k���P5��dslWS���y������z)�à`�'(tT�rn�T�4��kͱ����;��]�*0Qis[Wt��bC�>}�Pa�U����;�i��hgFf0�ӊ��g��{�Ҝ���.�د�[�Pi�M�v-K�͛��j���EG�$ʻ��V��h���OOk+iC͖�Q�ڬK�5��uv4)�����=i(��3L'�ò"$��I��.���u��2G��,�d���� J\��rY�V7aR������4�>�Ӭ.�J�/��A<����Wo�����	�cP�.~��3�b�	��z�y�ˏ�����iK=Jr�PG�"N��/&=Ò��վY�F�@��T��
~!x�i��Y��x�Ww�f:����R��X�Oi�F�A����6��"B�3�i7��!�>�i�mblTUS����Z�*?�s��S�p�49�ܼL��Rbis��������t���3��a����r�6�oP("2t��\������\9�٩V=꼜ڑ\/�%��{��
nI�xOk�1r2���Q�m�#����о���  o毑3Ӛ��0*�*#�Q�j���9g��2�+� ����]�G�}B���vo��[�l�!���v`���q'��-M���1�p�h8���y6�gY���F�l`�4{Z�W����-㭖8��_�'xW�}�	�ORlꁸ�)]U�,Uy6>�q>�hZ�8�Ҋ�Y2�4���|�b�jei������� ���uH�)��Q�Aҁ�sv�)�ƀ���a�����lz�A�F����n���
b����#�#�����z�̽K���%�����v�L?�'U�NK��Y�*���s���	��2�ղ�+���W9��Kg\�\�{���/�Ӥ�d��o<�w�tT��֙c��������KJSh�H�T5.o!m��ǟO��n�h��Q��u���d�1���_�_�s��k�h��H/��Z"��>ބkp�/�D�f��� �!ƒ��k1���t�	=�	�L �%{G����ϙ��ץ3�g���Y�~�ҫ�w���}!fR��8*z>C��l}J-��j6ʡ�l/�<;x Z��zb�Yh�TWE(c�,-(�.��>�����eB6����ڤ��͢w�͚��FdD��\�rRdP��(��sWK'Pn9�Q�O]~����xA���^5ܯ����z�?��E�����B0�;xA3�7�J�[�7��q+��bE>y�$+��ǯ���LT��~y��^�Y֮��^.!�՚��u�%K	��򒦗���V�:���$;�D<B]�w���`:���bQ[}�1�w ����Ͱ&��3>�(<��:���>9q]p��ށ���x��+�^y^�
�_a�u�����r>1o��s�ã�l/Y/��ÆRS_�P��=v��.T�S������tj��Ar|�}H ��:ޘw��6ͦw^ɢ.S��5B�QoB�SY���~��{���.�Vs>"�UgS��k����y�D����N�Y1��xB��I�>�|��!�=5NL�[�0#x$K{f�N�3K�X�U���hHص�&q�~\��u;m��׍{�ZÄi$h9�ʶ��}�;�A�\�ō��XC��c�uo���(������e�5 1M#�<I��*;�!��|�W���7#�	5f��l@����J�8*�&�`����y����Ő�~�w*�����`g��&�YWP�7���
NK|(��>/>x@�Vވ0��P�@��Y�r�����B�[����L��$�ﻍʬ�ǭ*�8���c��ܝ�G5Rs}��ݪ�.i�{û�@o�X�N���Ź �j^�p�^��IoXԞh��m�����n�?	ʋ�=�J(�fB=���K��p��ߏ0���%��%�w|6)�K�>3�F�-�s�Ö���Aasi�g�0ī�m ӌ�h�����4Hov�k���7�n�@<��;�>���M&Ed��G�������ˏI��w�FQ��ںg�B�z��[�W8i�K`�\�5��s٣$Q�#=�M�6�5�-C{��Xy����P��)s���:ӗBI4�o��[�;�����11���O�U����XQn�>��(O.��Ŋ����c"aR5�Zڟ�0�O���mDMmx �a�I
�
�S���*�'�J�0:J���A���t��`�(�r��{?���Q����h���o���c���Ĭҙ���!�����/��������Y�U�E����Z.߯���yd�ϋ�I�j[vҤ���h]��E��8e�f��L�
D����u�����C�c�f&d�^&����I9��mO�wt��TT�@��Q�������-YGw�~��s#�0�l���|t�fў��脼�����y܇�t5���7��IHLbX@�ټ[r�I��>��B��6�2@nWCoG	Yl��1�L���k*����ze�������mbq�ϡ��4�:�6�Z��6Μڃh�í³T�1W�V�ѱ, �E����:nQV�O����.�_J���:�y+���S� ��q���Ӹ�X��Twڡ�=���ѵK���HS}��眔�������b���O7����خq>/�`��M�X�K�b��X�w`����	m����F0�؍�e��zM�[��'$5J�X�~_�p��}�;�yD0�Wf�;�^B�]�Ǟ=�K�S�?�M#�pR���G���1@+GH���5qd��������[i����d� �J	�G�6�_���O��D+܍�^�����=?�E�1���F�W���y��}P�r���5�+�F�>���镯bE=b�WY�]W����ӯ����k����lF��${*���?:L}����L�R�(��j�R���y{�27AUOy
1��>�>$�j��<4��6�i���/��T-(�h��a��0��>��ךfNڅ-�(�4�1�o#[h�.�K��������^�6q���|+F��ʴ8�}~(�rD�A�Z!�'�nr��?P���UG��Y<.��E��c&|�>�K����a���z���������o��`ѷ�w��'/ �<���öJ!���txul/WG�$���AP�X1��t�_CP���B*'�y��q3���^X�@W����N4y��ʌ\�p�4z̇�ӸH��|Ӯ[�}hc�O�م��U-�y{Y�B���X��L^ߘ?�9���{Ƀz5�B��\��2HЗs0	���d�7�ㆆr�g`
�W8����&��dx��,�ʾ��D��(�Ƈij�(�~@9� �	�a~�@,��Gά��8���}k|##g�A�:!l�JN��Է�l�8X�&��3����\�-&)T���w\��@�5��<���҆o5|��v���M6��4&�z���|QӋGU��,��e?(st�DW[u��a�b�PP���Wt�GSӘ~�ۣ�$;��[Έ ��_��!���z���^�y�4�T���������(� K6��X���:��]lӸ�fa^D��С��ۈ�9��i-_;��v�����w˨��d�)y��S��{����t��?bA#g����OEZq��7���)i�}��׈�&7J��ϓ���5�@�~j)M����/3����4T[	�/���Y�A�i}f{�v���3��u��K9zZM��Ip��[�(p�����W��m"��W�cmO;i��Xs\�� F?i�WjkI��F�J�H$��
X�s�yg|x$q\�|2��&Q%v�;G�
��_�w+�����WcIӎ�<�$y-ۓ�(=kf�8��n�����㚣���b�=)�3~�ֳ���8���
cV_���� _�B���Q�
r���/Z�	�r@�Z,*�C��{@��B�UV|ן�+�=9�[F|��e��sX��qC���O�N�$-~���q�[1W>��%A�}}EEj?���
-Y[���{���E��� >+f2���D$�A���Í��$�-��t���דi�����#q��+�z�"BN�|������?��>L��/�6���G��KumZ�����g#34t4U�y4����Y�W��Y?ΣtV� ����;����ʊ*��d�������O�u^z:�ʭ���җ���N���VC�QX��8���ם�1[�d��N�a�ê��~�x��#����_qyZox	{�QT���q7�Y��g"�e%C!*�,�a��D/Ӓ�>h�#�G�3��]�%����j�\�=7�) �-de�3�L�T��?T�ct���
g&�Ll;s��5���ѱmLl���v&�m�vr:�������w׮]u�}�^��w
�����!;�"��Q�>��M��+GB�{�,>�p�~`LL����YaS���\g'm���-;�׹{���,����~\(����p"���eey����w�w�bF����Pu��ts�ZM=��6����G����GuZF�@=a'gԯ<�Y��4E�����2��W"FR#$4�#�ʟg:�R�v@�|�9��t����+YJ�.���wY������u��s��[��Ae�U6�0�
�������Z���{�H��i��V��h���'�CԚ����v�q�R{�����3�x����Ze��>�?u�|ez{��fBH��;4P�h/�Q_�_J�ﭛ֌�X�(b'���S�8[l#��P�rx�c%Me���,�&d�ؙ2~f��)�6FcB�q�P��2@WLS��́@y�ݗv]�k�����sH�90K�l#�����N�ۊ�k��l�M�@��V��W+65Et}[�X��zqn�31UϚW9�;%y<��y}6�g����e�G��I��I�  BA��ݵ>}��d!���.K�����T�wz��Ş��ܺYD�OR��8.Ш���a���(�r�8�P�z�,-	�8;(���3�W��&�_]%|J�����V�1i0�4"q�}��aA��E�-�a�'�w:�����1A��x�c����˝s�
�嬡C��;D2��e�����ߴ2�e��P jf�5-�tɞЭ^.?��vzh��R�T��l�>�d�1�(��M�	��9��s�]NP<X\/�{ܞZ�^Φ8�pq�1)��,`������r��\Yl�L�:4�M�k���|�];@���zq���`_eZ,��z�H	Qut*������VP�'�b�o�9<�ӑ��OE��<�;�Z��0����:niȑ�����g�b�ݘ������Q�Ö�yVt���3����M��[t��T�$�v]���Rܳ~|=�Uoh�%~�Y`���=TE ��
'����;��a��K�R�վ[ͶRx&?��#&d�3@p�G��H�8n��n����Ŝ�+�{�5=��g>����H��BC[��²n�\V��R��Y~V�߽�r9�̺ƿzu�"��xW��x�����7*2�^���c��}������W/��gr����m8���屆nu/ukS�"���'�� � r&ʕ�� �e�}�gXwϮ�� �n��d���p�^��O',��$<,�|�'3F�z?X��5�R��
���(�"uMH�aSSk��h���։��.��۱�u�&�ғ	�Sv3�?PQ�M�ޫq�1%��џw1��a-+������S1]��w􄈝�|�q!ࣷ��p��h�j����4���n��y���+?�J0@}�5���8ԆN��@����#��8{�j�>l����J)���)ڞe���E�n �|V(X �H(��GU@Y=:k��zu�(��^��9��j���t�w~��0�z7߱�q>O>$'J�W�	��C�eD�����T(f/-�2��}� ���s{ÖK|Xp,Р>)w� �x����ǩ��%�Ŵ���K�!JI&D��Y��f[
���<js����G���jbU�Z�_�?��-#I��k�y�Vu*����U��{�����z�=����<�� R�f�jҍY��Q�}����ҏYÍ��=�����[4�ˡqC*MP����p��{�3�y��C&*��B`�J� ���z��R�Wx=a�wU��*�_%�l��U6o�f�'��Ti:�u
�;�"�`�o�ٟY���ʷ��**6��Eh���j�ge��3�8-�M���^�r'�ȥ	���]*�2�'� �d6�`��y6}��VKHK�X�9�ϞI��@�Ӎ}x��4`������KA{S"�|�&��S�[R��g�NI�c	|un�\�<缵��?2^�-A�j��W��i+apS�($M����͘PXzMv��2N)K��uN�H��c5v@g�P*����� �!�!X���@��~��!�@mIH6���������7��?��b�����5��h�4��*����O�`���`�@Y���e)�E.�����wr�%/�P���4"Y���;��{gdq�ņ������X�A��ٳu��m�`�!v����+jN���v9��6����?*��
�K�����w��W3/M��(y�:2z��_��s���㙬2�ܼ���$����B��8�U/�֧����T�$���C(��j�B�	����S$Úor�@$�� �`��aT����p�X4%��=B��4��$���0�x�-dW��ɯT>8�V.k)����n�ګ��Q��Q��K�K^G)�����-2@"���c&�GD�j�|��3@�1��o�E���ܞ
�{k�Z��1Y\B~N[�X��3Ff���k*�(��K~]D���V�BH��{���'E㿔�=งW:���y�&���G��m�܉���O��A�3cc�A/ OHK�H)( Xr�sEsf�p�93��U�y�9��΄��w��o;8e@KK��t .�͂:�����OEB�y�VR�Z#�C��hT鷫�o�ڠ��s���C�M��n���R���Q��ߑ)7�mNЁ<p�s=3�3�6��C�bR৪�UW!rU<$;��W�P����o�V�no�gfS��ܸ	�:	;7d��L^+��C�|���r����4�KJJ�	��'2y��ѷn�u����~[X�
c�rQ�XZD�W�>�S<�wZ<y��/i,�� �N����z�����C��j�1���8�z�.N��~���%/�3***8�_��o/qiiaR�=V�;N�W.�J**
jj!����	?�p�O�b~�!�;��zx�rk|奭��9�)DT/�(V��q��������vjM�G�d��3,�R��곦1�8�L�Z�Mr=Wem�T�hR�	H���աĆ�S]�{����*��sZnCv�����A�X��V��Q]w�1v������ǌ���m����b��q�����P,T�Q(�YqJa�X�!@Dacά��&g��vZ��~ټ��H�j��V�-$�M�B��|m(�E�7�����O0����e���*(_�������pv���$A�׃� ˛���cvnN^UUTM���%)��yE61�v�
*�{�W�����Yl,�o�A�3���+��{ Fk-�\WGB?��=_�"�����{J������y7`��[������f����L�4	+kbI	�����ɝ��A��	W��8P!dʤ��
DQeeaII����'���w�5T����,�t�,H?Y�'hE������{O�̟E�PH����˩Ys�� sdw(.F���
h\���AO_1F�/�XI�����7���R����9�o`�M	c~��X��Tn?d9>k��RN%��g��PMy�.��<��_��%��%|�"GRy�Yy��u�;�ޚ��5@q3;;�=s48:*T���;�ɞ"5�����M`GGf�b�ݒa��EV��Z����;��g-$;�UE��tf�)_�_����UKF���0\4��+F���I���q11�W�x=������n}d
��x�n�x��	�z�A �)�k=o	���M��x����TΑs<q��֝fg(�.2�ʏ%���BI���c��������c
f�["C�?@�ofő�"��Ϩ���O�M�*+\")Ԭ��6h�JA)nY�l8B�\�kӛ�������v@A8�����#٬{�b�����1b�H\��;�6���o/N~KA�D���rY�Z�3D�Mn��K��H�F��x2�sG�
e�^)b!7����_+�N�Y3b\����k����b��1��8�v�P>�(�w7���QY"ʮ�$�����>��0�z����ъ�&W��<mN3ÞX,2��-�� h@�6�����.O�ž\}'m�D��Zˌ�rg:$F̗�H����(�נ�� d˯a� [�q �-����a�p�&A��v` ���!�i+1v�EK��אNИ3�{#�+�C*�'BuCaK�����N+��Ud�����y��B�C� Rl�E3콟C-��R��,���w$�Mk�e<�-/�Sf�Q�<�̜@�b�W�ϋ�JTy
Kڦ�7��U�u���TV3�r:B*�~gq����u���R��¿�>+ϙ3/�����V@AEu���L�'��y~��ȱhI�>V��ځ���#%�@���x(D�2֒�^���p_4),OD�-�R���s�3��B��t�]�<���'l���?�2,������I:��fୟ��esiC���b�8l��V�U��-�.F��̢��jX�8)���Yϳ,�{���Ι��T�I$��)_��1�t��k@׏Nl
������+f���n��TQ*J\�GP�9��!�ȕ&7��'�%��*t�l�3��-R5�1��^�����v�Tc��׺�M���'�aH���������&Ό���D�2s������n����=�\CJ��ؕ���U���?Y��[+�6p�-m�hI}�<,œ��{�A|n��tH@[�,�������J=|k���s͒Q7n߂~xwO4)M;
�`Hiw���j�z���#^+��Ȃ���R����ؖ�,*�Ir���W�φh��'���W.wTQ	��ȄVvXX�w����@�J��d�\=gy�m\6<6)˃J=R*R�A7�Zi|�eΘ
Z�2��Q9SU8w�?���$��,���#�8�!ݰH/{Ib��o6'؆�e_�I������U�abh[�>�\�0E�_F�SxW�b�
ݽdgQY�t#֟'���/���B��N(;���a�[��fN+M���̢�{ECH�Md1u��<=î|P��@�Y2c���&.�޺E�W]�$��-�&U�x@X�:�^�������_d��⯚A�E�*�.����UAGGGRrr}�4�V;�.]����߄���n���(o���3u�0�	���%��ǒ������g(h:�T4X�ŮP-oj(uʖ��T��9��ŗ��R�a-4y��h�R��8�l��7�>���)��H7^�=��������;�+�[��N}��.$����$�E���cň��ᄸ3�����{@1���SN��v�n$��V�B����U����2�pqS��4p��8V�ü2��6y��'b�T/Tf����ܾm�� E�E;ꝶ�p=,AT��X�0��p�GA�Ss���ӛc���[ç��fg*�S��#��%]-xfYl0f��#3�6�n�Q0+�&b����|�|�h�p��E��K+R5H��z2��,JFD�4pf^��U�fs'���s)��%��������Â7��%H��8��[Ai���a��)���L���XO�T�`��B��*�Bߘ5�:��'[�ƭ.��Z,�n���#!�a�3�΍���$�(���U��%�m��+��ec0��KX��s�Se�?�|�_\�sT�z'����M�hA�ķX#OLֿ!d}r\
�c�Ub�:Br�y=3TJ�ܮ��FG�ŵX�u�o�H�����G!IE�$���c�i p:J'�+�ɾq�V�V���b�o����Q1$��JG&���T��	��p�4���Q>��1O:Τ�t<����tqȵ1�OO�a��7�/S�2X5`*���8f���$?�`v��I��b���o�؞�!<5>�d[w���A�N�꒎~n�&�4�����͉�r0����7������`B�/�������o`�^|888U��FF�3�|�����,4�؁}�����xԌl
�ļ��i˧��b���My�(o,��t�5p�Ef�8�������Y@��%ew���A���9Ń���+9�k���qk� �����X�{���a�{N[�Y&w���H�ˑ���-?���Wdu�4#��,��cv�f:�w`z�]�i>�P��/Q�����2�՞9]@�LaoM"���B�ǻ�f�x!E���u+eqx(y������%H�����2N�4�������]�z�,ŝ�M�U�M,coc=H����V�q���6^XF&ajY	F��e�셁*�?�K��l�����\XEB�(�D ��X���l��S�GO�I.�i�ށ�g��F����&&҉Ͷ/�$�S��r ^[K6�q��^�*.�QT�m����4B��׭�Ž5��V}5 ��QSNO�-<��<ef�42#�ˋC/+(�v�8"$�}��;q��Y��F�4v�g�C�(PlCX�x�S��o3���³0�
�C~��4�
������
�t���Vy~��/�8<������tj"!L��%������	�󢺷l����m��|uݻy�<rx�
"�\^e�"%����~���U�]8�(o+��������aF�R}~W0��?h��X1��;���*�X3�Y��#����� �ϧNobC���r"L��܎1�ʮ'J좒�!(��ĸ��"(�	F���F�d�{�"��������p�mG�N�a��l'�R�rR��kWh��2���3�6yA12�E��'V�������׉�}#VJq�z���]�x"����?�f�/��@V��49����~ Z!U6�_���݀N�z�����Ys����_��z��o�J��-?�Iy5�硾����[��3�����I�ŀj���VM�"r������O������fF)T�X�,�k��%��෸�t_����K?FE9�hbc������/p�k��Т���s�_���~SC�(�0);᱐ݶ�R`B2��Μkf�b��g�ɛ�ճ�ж�!`a�. T�8b�M�I�wb�D\��.+Zzws����I0
m h�%��a�M���J?k�ʔ
y�8!�$� Rhu��IId��T��/�T5Ul��b�aA3&)��kƮC����^㔱�`�8�c�|�5Pf[8@-
I��X'.����C���bUk@b�d������Pr&&�/�寺w���AT[����WAU�;��k��J�����W���v��[��&�s,�$��`�����R�5��e��t�z|NO-L�d�̬���  Jπ'&-��L"��M0���Y�&r�,�B.!�� �ʉn�{ ��M��q6���L�5.���]�^����&��@[p����]���z��/mx�%���!K��ϸ�vP,�>,4���^�C55���]���ZW	[�g�A���A��^�*'7iZ�� ������,�L@�
�!��^��p3�C`��[�Iv�p
���i�%�]R6� ��q�`����DC(��3��O�o2Җ������fl��*�b�m
è�	��o{�!퉡�Rv��hgQ)I UR1���pTV:���P2�������^K���0�Td���e.דomxvX��Ic�X�N.��D�R�U�/2�^�o�^H�X��5�STtEL'n����WE��+۬�RX�M��M_f��)�$G���FM�S,�9�wve���S��wG�@��,�ϧ��J��3�I�Y���_�6��6��2�ph���9�o�c�G�B���?[�4lЃ�����Isy�����v�(�ϦS���CD���r��
�2��נ�0����/1���6/��wG�
������z�M�P3���TZ�N@�C��ƅ{4�|g ��H��А����n��t�Œ�E����yr�hM�Ӓ��^U���/�26J�	��@v��'o��E�JY�����O��
�"�&���ZR�=��'�f&?zr�2a#�IJQ�W��Y���j@rH���WM�2|(Z�����ǧ��>2���Hތ��n�g!^Z�uP�b3��b�F�q!���A]!��/�y��\��?��(�0�
ʞy��ǱyK�: ��� �{b�H�r,HPj�Mr�%���sj�T"��o�5����g'#���\v,�Z��< ��(�n��[R�vQ1�O}n#�:��?Y��mJHjA.8{_�����MaR2���6"���wN��,e�F�0>%E��b��m+�������b���c8�	8K���_jI�!�n0�p�3��|jMPʔ3�
mm�R�0[��lQ��CʋӐ7���98��qc��H�_�e�c�� �Z3�GPn�(�?�b�G0(�\��
$�V�
���6`c�dY��D)�%\�J8@\�� ���D�k?�2�X��9���"
����|��t&S�a���hZ�X��g�'��N>��>� ��7o����x��s'�p�}��,6�S���1�ߟn�e�'k�/�"V�k�g��.̏��K�P�7�G�Y����nrE���d��Y+'�J��T�����X2�M���Η(=ۋM,tQ��݁6P��gO�-��X�{�Y� Գ}��b
\ �pL��aj!XV����;��"���w��{/�����|+5��둝ʂ5>@�"�bC�3Z:~�pF2SGhL5�t�ǟJrS�+A��/p���I����`�qa�f&P#�v˅���čQ;�.ݵğ8��*�H\褡�0��殚B�����>���jxq�iG
�pq4g(W=n�W";7qз3�C	7��SO^2�OV|��T{'f�D-{Hzz�x��z���WZ�`��#��p;k1���.c1h��0ľJk����$P��*⌓����S��Ye{���{n�j�F?R��Q~[5�I�;����0���ijj=d08:�/�w�A���3�7�Ncrr�Z���@k�Έ(��Z�_�r����KbqD�]�l�P�?�.t1rYaˡ'uP��T�4��s�_.�L�7a��67���J�.]Nt��U.�_H��VQ�6Z�CM��Z2����}@k�b�(.��m��򚭜n������+9=�Q��̐`�����+��БiY=#O���vr�i��f�Z�~��]s���.Q�Wb?$�.H��X0@P��XݠѶײ��{�h��f`���TX�ڜ�U�贚�M��6M���<�t�hR]���*iV���7���,"$7�8��S�f�!_�aϱ�`'u��0�e�0���|��/�M��_'!G��zѼN}\�`�Դ���C�p��H��a�a��2 u�Q�QQp�/W������_�uE�r���^-��[��w�f�T� ���6������������^�jOT �~�Ja��l<ޛf݁]{�t@�A�"�h��4�-^5F����A^���8��6����!J� ���f�)[����3�:��VE'�<�����7�ۮY�l�g*iF��/c�x&�ᏼ-$��cxhO9~F���w���_|4�f�$�p���1T�[���_b��7D���?�G�&�_-	R����~�:�T�����r=�5qN +K䔵�{iMo�-��T���I�(P�6@e{�|D+T,ea/S�^u��I�B؋aT�Vr�ƍ̈�������w����o��M�z|�=���/�ڀ�5J��a�w;�f�x�xs
�,d�ha�ɰ'�~����O�WFZmW�wFd>�NJ���
��Q0~H9Rm��Q��_lwc�%6�%�����\��r�߻�q�ɤ�X��b!��ъ]&��"��}��^���Ťx� \�A{�q��v��a̳AG���`Wbi�ѼIndK+P���t ��Uz@����	��N��GJƮ"&�(�-�Llƌπ,_T]<�փ&�<v�'x�R�-�ڿBķ'
��	Ʉ�&�A����S��R>msػ>3�S!VN߼����C;�U�)�o�;Z>�	R�:��90`xD�{�0�@K�e��x�X����b�a-�����+��8��V���4�~�����lY�O@���$��qZ�]k����A��ct�h��c�bB+c�5���Ci�s�#J�A?�d�8�r�D�������<��an��?��9��_z��'�90�H�c2���R�d�E��x�w@�ǳ� 1gՃY]�����vik?�.�\dG�,kF��J��"�%���؀B�!9N��ޅ 5�1���m�4�ؐ$rP�-B)4�)�j��Z�4��[����h��s����
H-P��%��#��}����E	�p��f
󪪐�` =���,6:�s�T�ѭ:ߜ<@���9q{8?�%���ot9É�lr������3f��e�%��o�7J������@�Ey���b,G"Pr���Y=��l�?<I��󬬷_�0��K8!�A0,?C�i���_�(���-˿F��--f�6힐��Mǩ���3���q&�`T�+����)����ewǾ�@���@Cwن��2O�ӜkZ����246�˧��8�Q�`i ��5�XU��Y�퇨e%1����TVQc�*�u]����ڹ�q{��W��;��	�^��U�K��:s���r�0Oī��54wN	��^�[Oo��#��e�v�R��>��QN��%=���s~M9:�B��Ke�x��KjG>j��V@vݫN"7,��E�M�/D/��q�~J�I���)?  @��!��i,^��B���X�s�Y�I�j�̦��/QE��\M_���B�A�X�a`B��Iv�.�*�.RW'16ͯ��Ve0w�U4�Rͮ5���1�5���Ec�vN^ZR�c[���'���t��ja�jY�f0樦�ry4�j �	���9�T�XB2k.�Tp��-A{b�[g����	����|�q�R��^1�,�����"j�P�~̇�ګl���h|����j��f��Zo"���9��<#�͗�#�Iq��N��'SM/���v�'�~�R��NX����M��)�1���S~5\9�A�\�5�Hk�/�K8��1����w�E<n)�ܵ߂��>��D��c��n��G�:�ڈ��R.�������k�yT�5�T	�7����B�y����1[���|y'�xNPe-���揵9xY3��<'�UK���晛�-�V'�� k��>�H�����اR��;�3��ƗS̺|�;�}�#��m~uE�ry��xP�_�H����u8����Af�_�鋒�b��罧���1 b%հ2�Gte�Ԍ�Qx9�h�#�I�,� R��Zi�؋$ڌ��(��v8���.����;:�jQ�%�X�՚��.����N�E�|Mr�ͩ�ir��������N���Z
�g�������EL��4�N�i���D<+Y"��M���ȝHY��C��ѓ_�ʒ	H%֨S�( 7����e��8�n�Vv_�l߼3�话�-�7���UR 4�m��/�ٍ���)2�
�lf8�U�����j8MJ�����Ɩ�T
��ݡ8��?U�F ��Zu�j��6lG�3a1Ș¢����L��i6��l%�@�YU��CK�#� J��A*�ꯁ��}�@=˳/�H��A������-��]���=_��Q�Ha/0�6xI))"��ڤ�"q��(��Y�߹���N=G���$�d�"]3y��/"b���l �)2L��(�E�ɋ"A�q�	�jv��Y�=4aE(�ڿn��B�0�p�(ǻi�:O[�
ӧ���0:qk��'�/�8p�.�<�|g��F�´=l��$�Q�{B��n%j��͊n9_s/�{����U�C*�Y���!v^R�[C<3�"C�M+l6��[����� �����ΝwH	��ӢI�pS�lp�u���*j�d\��c���U.n�2�������I,��w�}Z8�����I���ɻ�A񡵈4�U@b����&�JU���2/[Y�m{�r�m���B�?NP~G������z��c�֜%�"�%E΀L���p��C��5�K����עR)��?u,��'e�nw������.�o��fM#"5�˿k��Y�N!�ރ�>=^YC3'��J}���k|���(��ĵ�VQ�R�@��Z�Z1�V�-����F���Aae��9M¾y#9x!�C���=�U������۹�8�1Nrb�W�+�Y�t�{�w[`�z_��{�I|V�����纈�`vw�9��x��Ͳ�R���IM��(Y��I�˱�cHh:�-��%z����J�׬�0�����mþ�8u�h�"8�T��F,!�H���n���"B���x���u��a;׹U@��
�Ȃz+D�l8�U�#i*�Aע6�ȖT�̯�5�In�6+	t	�/A�����aW�G�kT[�E�9.�15���,�9Qq�}ԺMm��t:N����X�OI�X�0W���|X�3}�Z�VK�GE�rO�[��1����q\���öj��#�_(��f@��H�s���^3���r�3Ca����y���\
���:�}:w�Ĕ�T���h>�E1�iP%% pJ�s��=m}��q��y��wR2vt��]^G��\��ux%���+�p����[��v���V��M���_��zū�U~��R26p���='�]z���7��n�|' ˚UW�h�MO�ylVSSc��miIG���������������A�W{��˹�$�Xjg7��͗�����nB�ӷ���rg>.#��S�\��0	ژ�u�g�r�D�n�gmH�?.��r���;��t��S�:�ݍ���|�k(���f?����R �Ht1�^���K���0U>Y�mϱ�d.��<fVʪ�٫Bu�+���V
��.��1vXOg�SVV��0ӹiʮ�itFud9ﯙ��Y�j0�p�U�i���3�m�,�h-EC�VW �ܳ�lN�P]��<����I�:���8{�'�\���
u�i�<��@լ�(?�(lP���%�U�P��M=��O�w-~�������Պ�%�C��pB�X�����i�B�`u�'�4��N��=�3A��-��[�\�ٞ���ϰ`S���Oȸo%6
c�R7'�#7U�4[��m�p}�ƭk蟨�OFZw꾬u���
��!��: Q5p�r�����a}�ɳ�S<z�7�?��I��L
P:[vHJ���Ek"��'W�G�'PJudp�c�]e��*ng�@A�˶`H��P����}�z�I��m�~�3��.h54,���?0�8 *=%̢�>���r�'�+s?�P���*a��7U��p��I��;��D�t��:��]	r��#����+��zZK=��b?zo�A8�����`��@s�����L�?��
�G�A�@���fϤ|>�ͣ��	�ч�j�JdE�L�W�C����F�<ںfr�i�/�w<%H�ᒁK!;=^���u?��ϣ03V��\�s�o����m��ey4�@��� ��u�*g��z�q�O�>�jR�i ?�YϏ?��2R;[.��o�9S�d���N�ɜ��ra�;���c�5��R~�:�b]0�x�
%�fR��w��6쌗oT�Qr��j�������C!t�C��ۙ���)!��I�w�Vc�z��&�<돆����Mk��$?���ܪj�Z�~/Q�Z�ױ�Mg=W��}�����V�j��Al�}Y���x�շ�����6�h�=}���<O�c�Nn���H�\�U�6t�\�Ql��r�ܢ�~���z<�+�9cV�.{���j`)+pi��D��o�>�N��6�n�ˇM�͝�'C��d�#���w#w�#Lc�c�F+x���:�O����U)auhS��YBz�63����Ǡ��nO�C�#%z����$����2�Ձ�tp쇉�7r��:��q�0�pV���>1�S�E���D	�_��p�۲UZ�����b{L(���Eܪ����v	 ���zo{U <[춆	q�	n(ӾI˫Vf��IΝS���xil��6L/��kj�i��
�-BF���8�JX�J��؍�ll,�\����n
�7x�|g���9l����uV(G�*H|��ja�|�=�/w��]��U���}	�Az���Q�=]�+�Oˉ?�����~��Wի�e��:~�cyLLG�-� �����2%\�2����q��]C���s\�~'��q��:+�#�.f8�DB�.I�K��.i��o�ޞ��p��2u�3��G�D�������k����Yr3����X�/�fRԞ;�|��5�2�^ofW�<w�S�Q�f�ڟ6Ѿ�)��SN��q]���N>~ڬd/g9.��������G=�sp���ѳ���d��Ӑ�����*����H��� X�ϸ��#+?���W��q.o�B�V��Y��QQ��B���C2���2��4ʵ�������Dt4������P�h�S���M-�L�W����ﮰ�iݒ/T��<�j4� ?�
��S���G�i+��^.�˅�:ϻJ�P���o�t��_������Oˇ��2�e�
�,�"���I�2W"=�?'�K�F�*�KBgn�������Kf�@�����t�Q���"�r~��ig�8�m�.;^F�����w�ZE�w�˴�tpMq��98���A|fe-�[3�I�Fi��NK����$�29���ĖR��d-�d��n��6�� ,@����ֿ�G8>����/��_5����\\�r����JVr�)�~
�:��W��I�Bn������	�rJ�֪/���Jf��jJ����Q�oe��.�p����gR6
1�d���e�9I��$�s��?��aO�e�cQ�����~�����X2�=9��/�33$-Q:(AWS��[�9�M'��Eʹ���^4���͗v�D��)h0�9��S ��A��TݭQ�D�p���}�k��9g��w��i��H��0f�O(K�	t]�K���R�p
����$O�*	��!7�8W��hT �.��ָ�]dmsO�z��O���	�)jch����#��{�/1��rZt#��|=꣭/�v��� �v���'�y�f0��E3�4��݂bMBp��bvsw1J�����kb[}k��;�_����� �¦�n�*�⨝HJc��.�*��aG�E���R�h%;��M�h���oA�p���V���N�k�p���I�
��(�kr�Y)�W#H�i��\
�w�� a�mM.�)�!�ʔ�A?|WO2��W���i�Z
��߇ҿ?����6^XȤH�
#�u��\�Q�$��i���d�K�t����D�܈��Y��(2^#�Lb�8�*|�����u��z��8���%R�U�zÊ��&�$f�[eSē�L��ە���k����Y0<��t�_��|�x7��3�C��+i���x�w)5�|���}�L�����ܸi_�0�,��oUy�C���9�A��t���0q�E]��<X��W�{�-�2��/� xT�^anrB��]��~�,�a�#�З(P1?�Q=�p�E&ԏ"#��Xe���r�-$$���Ǹp�O�d���a��ݺU���l�M��c�w�H� ,�K��fU-�߶�Hx*u�*�kB�T�U�9���C��6��R�����n���ֵ����(Hf~G�xT6A V�L{����U�xO��{���6e���U��>/+�����t��o��#S�J����j�
5e�\��hWb�̗zz�H��UXSMB��i�^V	{+����u��-���!��.�Ҏd��ɍ΅�2�Q�7O$K�u2rgS�P�{Q�Y�0�ʒ6�����%fi�t��,�+�!O
�WE�����q���G�K!��*4#�*��/�gKUF[�@:�oV����S�mJ�+���c:m�Y�\�BO/��א�X�%�"����9v͢�kC��2�8�gR��r�)Z�û��F{�j��ٌ�ߌK1��:��f�u��˒eT9�)I*w<˩-=��A�{��S%5P��zx��.)�L����a����b��hu�B�h�e��X�9P���9�}�Z�"{�4��
�F�flB�j�k��<��D츍��o�E��vz SI;��d��h�|���ל�f�l���G� �7��A��_�%=?hҏ�3��=^�H�y�}��s�r}w���}���5���ݶ����mp�Quʽn;�Y�`r�p��Ѝl��!�cGz�������!`ĭpmE��
�#��a��=��(�Qw	��<��k�� nu6���J�#�%>ʇ��y�g9�~|��1C��P�V/Q(T�_y��V󥖌�����`��2�?L
m����Bܰ:��&��d)�w^���4�ANp�Ḱ��-_����OǷ��_U�~�복b���jM�p&�����|rAj��w���}S@�c�LX�-����/ɬ�hi'5�6���8���t�p�j����EHX�V�2d���u���z~D�Ь��9hP%����G�Ðf,������L���_.`��S��yS�8$���{��^��{=��][��:��v�1�U�pL���v媷��kUYw�����h��BFF�Eݚ�,�-���> ��r�-}��-��:��J�2�E��09k}�5�-R���c��=hl��d{"R�B��~u�1`2�W*O�F�w$+ӾkE�A鯣��P���Z�h��b�#D����/-9���qh�D��bW�)���Y�t��Ll;�ض3�v&v2AǶm�v&�m[_��w�?�G�}v�}�VU�uz_�.=����/Byr��z�e�鈿�GX2M�C�-3h��Y��U��<�
���a|�d�C�N�[�a4�ԙ�%��'xP(c�'��a�c�j��R�����W���]#�#R՛aڬ0[h-��"M�e�t�֜
��,�znd������I稦��q���X���@��=v�9�q��ɻ�®�#n�"�0=c��d4jU�!g����4����|+����u��v�;���hi
�p����f�� .rY\Ǻ���p�@�d�Ɣ9���^��Kゐz���+���ۿ���[Ƥ.�
뢌鬍Q�	M�I�?���	��n��536�(@&�+�|��ٗ�f���`>0 ���K�N���_8�,ۄ��~CpmE�loa�t'�ܞG�����U��L!������"�E�m�o����%��ѳ������	��-]`���~������r"�zg���yo?�ʝo�ȷ���M��ۍ��[�Cp������ڶ��Vʅ���9q�x�H�*7n��o��̈F}h�ß������&S4&,C�w�b�*+��' �̵[��(b0���?l������+��q�f5��_Hc�QWꈃ.�1/v��Q�,O ��R�^3�`:��Mh���1�f8�`9+��;W+��=5#�9~����F�=�ˌ�"iK�)%.�/��Ϩ��0'��Ec2$;u�ޣ��,���M�p�*7��v�@0�E����E�	��v4���<#F�d�p�0���uE;%�>�b�Z%�f�c3c�a"�6ϣ2�n��4�~�R�ƿ���P�N�T,k��3��Cp����*~���`���b��Gj�Үd��r��q{a�W_�X��&u��\�w���o���#��iƭp,���	�ab�z��<ц��h��}.���)�Ov8/m���r�O=�OR�tiD-�X�Kͧ�]���r�B��fJ�t����@����Z�	�*31>!N67�/qee �,�"���;۷�y�퇯�e�����ᷲv�z�B�+�{�'�������|��(��4���
�ƾ��t��s�ա�Ԗ��Z<E3�}2R���-���|zT���$��K8;;;��=���64$A����%�B��F3ϫ2�F5ș!a$o�L�"B����&��֊���An�|N����z�9C��|)�׾��|���洅�`U[u�R[����������Y޺��q0N��c�3 �)xGy�=�&_|ЁI�9�TY,"y�M;)��,�h��ttq�����v+�i-%/�g��A�XH��R�c�����p��-u�,�����g�L4sD	�8) ى��Q�W�w��[< ��H�=	$7��9��^i[�u�8�x�{��|O��7e�0�#�{8����=j�fz���GTɠ!3��rx�FX.p��ʮ���3�)Wx��l�Y�Z)�3���m���r���˥[������3��Ե��ujw���J��=�Y�VHk��t�ٝ�6w{m���o�?�p��CT��ZJ�풤��a֙��(V����`v�R�̄����b��]2������HY�Ʈ�K"���i�))JV��������-ʂ��Z�-�.�W�D#�i�J{���-��t��b��qi�U�H����JI7�'Q�<w�_��JWo^���	JU�a��ʷ���8mz�!|�*��:��}�7�� ���@}[j*x�r@����n�ㆅl�Մ
F�:+P	pox�����gi���{8W�0�P�Z ��A���FW	�`�m'�h�4iŵJ{���	{�.Z O{�vn)��ݫ��	����e,�R��
�@����A1n��}ؼCpm��Q�`�2����bQ%y	�qP!E�]�	�x
�叮Vy�Ѻ|�%Ѿ>��T(o��e<*B����x��NM20+	����:L���I1�x��H`"c|j?�̣�W�ͷ�%
$�+�n$%&��n5|��Ն5��02�n�؍��}��k�F��S�����G�8�� ���|�Q5����Sƕ6�-ڝ�뷅.lt_4��ς��<z���ڪ�#�
���q�j��P�E����gP/���s�2CJ�!�r����ѥ���:����J�M9���Q$�8�:53T *|�gU�:���nJ����-Z~�P����->γ����t`������fG+�"̰�V�A�A+�bR��+���k�3��O(4Z>�h���f���J��y���HM+��a`���C���F�V���]
��
ƽ�w�UI4��vo ��lk�Կ `+D@9��F��X:C�N|����u�}��!��~�SG�&JFV�\ &�1� ��Qw0~1���)`߱q���C�7���r���n�A����ﲉ�-.r�}�ږ�]�IՃ�#�nH�)���g���7�}-0�Y�l.���+ش��G8C%�6ZD��sJ�-G�a���B���S-/S~1�k�3zj~X��-�#��.���E�:Y~L�g�rI7�-�\���j���������}Pf2���_�Z�Q\e���h�Z��ͳ�)�Ȭ~s>��fݡ
�H�?�ˣ�{p�<^QZe�52�����I���5�ߧh��M�$��N��$�U/�����@
5̺��1�
]�hN���0������=��� ��c�!�n,eݽ����m�b���,0�J��n��9�x�����"?��&Dhv�#���g{�����
�����)�����s��&�
�ߊ�v������ׇZx���EeT����K2��(��o3Ӂ\!����L�G����߫p�pJ���zJK�^��#�~�:�/�����S��=������;�&��O@=[/d���T蔬lh��lW^����w�<�ir�IV�>'��ཱྀ1�2�sg�w0!��CC�o����4�ۚ���0��.@u�`��m`�,������q��\b{C⮽-Y����!o��Nܘ�`��a&���C��4뫃�!8�ô�Ba���Kˆ���)^k���y��s�����2/Nd�`�_5��j�IZ`��F(�1��H��1�-�=��>�(>?h5��!�a��c��6��q��h�p�'�m	"َ-�����R�B(��v����Dc�7\m1�#~�f���z��xcK_�p���`���t�-v,M,镗��}K\��[��l���w�ۄ\J��ݚ�n8ї���H�Rի䎭P��LB�KA�<��QwM�^M$Ω�Edv�����]5۴�@~��$Y׃�8~t�����Ҳ�J���aw�ɛ6�Z����!��Q��+w�"����
�e����P�fX��AR��
"��~��D_}��l�ڍn�*r�":T]���e��@���/�~ ��9�P҃�^q3�~A߁�n�dv��X��3���pa�$;<���:�IǺ������wy_�T2b��\&%XF���"t0p
:�_�_�U��OS�"��sW��F��X�]7�phO��۵�a��;@B���Gr��4+N�����3���)�^a��޸K��i.+�*�1l���ʌ�I���xgb�ېv��̍�	�`�u�����������P#��M�ӵ����B�o�������Ir����ی)�)7;񥱤0�����,v�	��?K�& 1�ϥb���l���ų}dk*�@�zM�ǹ�i/�y�(�o�����Y�\�WH��	1j%��^&�o+�ܵ���ˁw���V���X>X�����Z�>D���x�ҳT�+ti$p��w����r`����:��B�����"�����S���S,D������ֵ�'3lW6U��(�="Y��7ҥ�F�a�U?8�����	i����C$�hy'!�����:D��^T/� W�"�=��	S6+E��A�ڄl[�ad����'�� �A��]��1�*sr�ݧ�5��e���I)���!P�W�������x����`Ō���p��,�1����x@7/vn�7e;��VQ�m�@9�%L
+��8�m
6W���j�`�����!�P�V^���ܒl4𚥳�WA��[���������@^O�A�<���s�G��]S����?%mv]�I�9�r19,��X�vG���g'.�|O��:m��F1�W�kǣ(@!̋YP�Z�S��e��������<�4��HuXn������@�W�@A���&�s~��a�4�Q���-M@�z)7�D��LN4�r�So�b�	33���z���w�`�F���v���M�����g�yï��ˑLBk����g�d����P�b!�{~%:��*#�r���Q:��/��Yέ�;�'�∻��nq����Ol���^�&O�^q��{�-�h�� @Y��tr6rG��~u ����)�$n�0L!��OL+���(�,
u����
;��M���L�a��v�JڴT�޺�1��S;-F�Jw�K��3!a��O�X)�w���<#���D��Q�Gw��L��jW�E��vK���i�j��ޝ:�`WKŠ�aUj�C�����Xk����j�?�J|wOڸS�۠�E�z�%��^8�JP���J���/R�Iq ���x�,���M �Շ��E�]|LrT�NG�S��2�����(���B� v�8���'�<E��^��97nm��CF#�ex��'4��Zj��^�G��iFψF��R�\^�I�C����i�^a�m\�(� xᢻ:�}/����V�E��V�� ��ۺ�d���j�����DH��/��_�/���8��嚬�8�;���^��'�y����݊��i��Ĕ�MD\iথ�8{�U\W��u�bg1'y��k[�@���t�����-R��wD�s'T�|�=�q� \x����~ֶ,z7��ɜn�5�!��D�����vd�ۘũF��?2�EVV�O���쪋0 �E:�@2P���A�2�/���=K~Dz�2��h�����<-V7��ªU�Ere������$��:�v3ch��]�.�J ��h�P0F_1���b|X�>2�l�8����:����K&O��ѿ��%[H���J�aI��W�y����2���J�HFO�X�Ÿ��ȧw{i�M,8IA&�F�U�3J�ecZ��a�uӂ$�*o�"�U����4��O�����(Q�� �dt���K�f�����{���{���G7v���h�HM�;��m���*Wyn���ZH��;��n�W��_�mJoJ���p�!$Xh��@t�pw	Y��5b�pU$|�)���ۏ����A�C�h�*���37�zը����9�sC_��K�x�!��5�\����s���������ǯ��0���Q����˲*+��Ktt��[�������:��R��sČ�������:���d��Q����R,S6t�?x�#�×U�8�Vu\��49����`���D���T螩m���՘��Ҵ�g1�ǩ�	)�`�zYes��/�?�X���)?B	��M������$��Zs���k)]E��gX)�M���QN^��KjZ�E|mM����>��3N]c}����cBa�A�T�V�Xn�*c8ȹ��
r����o����m��Zu�y$�g���7Q�4_u����!|Tk�Nͩ�7��89�r, '��*�)�0:��@��D%K��STCR�Қw_hм��m'��2��� ��}��7��N:�D�d��x�������o��<��؄��K2�V3������K��]S��F�8���?�W�I�B�XǗR)"|�Rp��'�y���(.�'Alҋl\'N�.��36��+v��@v�1s�Q��x���Ee
�;}���pc	}0�#���<�E���;"/ޢ�I]�!;
1K�f�7���RP"- ҆���U�17��Y����'�J�Ɯ�y삵�(�󞬃���##��XY��ꫦ�*�뙘��Y�y(^��'�x�a�����aZM��M�  ��6x��1HRwF3�Z��q�УQ��)�t�yz��5F��[t�> ������8��L�陛�9���36��4���}�a��(�g(a��M>EA�I��c�W�����7SIi-���p�S�w�f���.�����Y�వ�D�BX��q[�SwC;��r��_�)p�j�je}ԝ��ER�|��qXnL�,�΢��|�^��ܰ�+{��KG)])��~���N#�\�c8�!���FLDI�t	K5�Y��$ozw9�y���/~�qx�K��B�L���"*�����&��~�Br��W<����rTi��h�E���0�f�;k���;����-��k�f'�5��,}S��u�KR�.�)���m��`�OU�9e6�;1���(W�H��^HQ"�ĩ/�i+�q���B(R�X�?��6�~-�EX�J9�}j�j�W�M�Z�֥p��t|�*�� s��P�^rI�n����ԯ$/�bV[�����D@
��Iml�gR.8Ƶ��c�, 3�өq>�LU���<FLs�N���ځ��DX��ɠ^���O 8_�YP���!�Ե$���w��	�X�$C�iDv�q�̹�����gfؘ���RR�EG�63�[OK�a@�F��	 ������cǘ{Nv��LݮW&wz�M�(�d�
JO��zؚ�2 �@Jo���$; �ho����R�$\A���E��S�L���Ƃڶ5̊P��W93�^!p|"�(̤�Q��-�P��>��wg�2�rM(�}�6[�3�챩��$�k����OM���}�R6,4���N��#�9�-f�w��RBIR�'<�������m�5?�U7������3[�?�f���}sښU/].��G��d��)^׻�;	��{Q� �P����,���_ƴ|<P��6��{'df��7�ɩ �	?��ʅ��!�������bJTz�M��6� ���S��L���}�B�pdz\��.Z6�d���'ڄ��No��"��M��HAҖ|X����U�FL9�_��_��<�kކ*Jn%3�E���-sX�g)���i�!zAR��\�s�=P���ձb����
j)�8k��h-㥍,	n�����Ee�}���#���!!�����,�%�Lq���m�n+W\�wp�z·#�y�U�����9�MO�B�X]��^����3��xMA2�(��63Y�~�_q7ҘS��$8�q �����]>UE�!!��t7`q�<\PՓ)��ꦘ�@W�A���g�'��e�۽�5��۰{�-��%����Ի�d>ջ�E���W{��z���3.��D- �fJ�O�+��&�I�w�s�K�?�����y\=�Eрv���Τ��������\�Fm�c �a6�.	�(~]�9��Q�$��p��;~������Asq<�H��h�}����$B{�¦��G�R�"�6��&��2���޹p
t�@\�B6ՋN*�~e�8�{��Z�U�y���o����􇒲rlb�7�j����&)i���L�*;�r�l�T|q��T�k㔛_�ʣ����p��yj%�G���,�+�~�ܜD��e4G�IH��7ٟb�a�;���<��Y��~���_j����D�{�¡�5�ރ�j+�D
�V�J/�?)k�,E���+��*�����������\L vǶ��4�܏	��VMi`������r�I�7-��25J%\����1hQL�a�3;Z�����hic!x����4K��>n��4@!���	]��8C]釄�t�
b޵�C��7p?Z��q��l�M�u�����C>l�������x����m�]�p/������8Pʅ�{����EI1��(��ә��n=�}j,@�A��@*_Nl}���ۯ�q��ld�F��`�o�K��P����6ͭ(���[��Q#�����}�xy�N-ߦ37��D����	�����R��$�/d���$7�DD`�P=��␉��/���5�����:��>�1G��[Y���8������[]��3<�V��'W,��dKmbEc���ݮD��(*;/\)�4��~��8Rp�RL����T��|3n��p��w�o�c7r�T)��5K��]��d�QB���y�J����滵%�D�y��֧iٴ�$�=T2z��Z񀱶1�
j���w�KA����멭�Nm���8d�'���� %k�Z�������ͳ��r[���gq�(����X�h1��8u&u�����[�Z�7U��[���U���	S>۳q:UE��p+):߮�"(��6Q���z�u��RI��eM"vwu_�_���2��gjJFn
#�$[���5�T�b�/�Lh�����>F?��&��.��B[J��f)��M�ԕ2�$����O�\�g��\f	z�x)  W=M��S!Q���`-����'��wY�'8%�%E�L4>�JvC�d�$O��!�o�J�����\\H��\3]���	���d���J��5B')�^~��[�����P7��==��+p=|hF�:��}E$�J	�(���H$O��Z�k�W_{�{�}Ĳ�T*5
�1J�=�h�HB� ���12|��m��{/n��POz��ǵ�i�FѰ��WK�@
lJ_F��~�-��`�d��� a����c��(Z�)�/����5�צVj��7 :�{baӥ�������QY����Ma7zF��.�+#�l�N��TrfL�Ж���w֖�V����0�?aW:����Ά�lo��=a���F����j�}�ۢ<����a��GS�0kc��s�0M��v~-�T�V� �fU������Ⱦw��h����+9ƍIO�D��0��`J2f͞�r��
��YG�ž���C�����7l5)��׊�db��X/�PB�o `�~������e*�[����1��Z[��X;�NM�:6<�����<bu3_�4�Z�Kl��c�A4��l���m�˻�m���S
!��]9?��Cj%�\W��{����Z��vU��g��`�"W!F���JW���!��X�zI�r���]�ˊ]S���k��T�K��A��Z͝����]¤(Ojm��a���'ٓ�ᰳ%���~-դe�8��Ԥ����!T���h+���|8;��&P��^.t(�e�B� :Q9�S������I�Q�������U�9�Sܜ��Ƶ���RB� �	�+0�W^�
��'Wd����(3X���o����[�*V��c������s7�Ra�R>��y�;�{g>�_VR2��0�k?*X���{���U1�e�n���v���n��?�%�U�Ĥ��y<|�?^*`܀�E�1}��mι��ʤr9�Vʟ��ww�)�9�d�yqi
��_s����@j��3����:^ж�,�R΂?�r�����AC9 [G%�J\~���ܺ��ʣ͸)���D��Y�xK�9��k�ń4���z�ll��Շ%��9���
c.x��,o�����i��т���?�O(�����P4�Y��zz��h��4��
�T1	n�.���o�~�#!EB�4��9�T?
�O�`lW��t�B��Y~��ԕ22�������w����I��s�7Dm�l�z��"Q��VU�\NkQ����jU�u#��������b���cҸ�`�U{q�2��x�`n'�RLʉU[�	�9�1f�Ul�Hd����������L2\�.�n�[����I��`K�_�d/�2"u�h�^���� '�shd_x��u��}LƤ"H�@�viʡ��α��+KS�xf��eI�,���I��keͨBS����e�*���-�RMهr1�;�����H�Q��I,�x�z�.ʢZ]�].�UZ
�(��~&j�\�;�!%�*�a ����y�ۢ#N��	�g�,�S��w2D�JͬЫ~�<QJ�#���5n#�]T��Z�I�;�ǿ�:o�,�}k;*���`�Җ$O�|v6���t�G`������m�bA�S4�v\_P��Vy;ѧw���Vj�E���k8�]EoYk��\Cl-O~��TU#"q�1�2�L�yرJ�T�<:�R���W�~R@��f���5�����q��"�$����w�tow���ZS���z�@e�Re���޿��K�i�Im�Q&��Fxu'������u�F(���z/�"}�!�hA����?����笮"PRxw��W�2'i�8�5M�)��z�}�W$�^v�p���4�J�U�����0Wf�24���PK)�G�If��e�4��Lþ�eJ�zvti���[`v�K;�U�� ���jU��[=)⧗�g�WH�q��k.�a�c�'�V����`��?#Cִ�'$j�Q��k1
Q-;��t;����s�H1��;��
5���E�5�.#˩��(;�> O���q���a��Hv=e���I�Χꨖۿ�
�T��u.��MZ$�q�':"��YӚ�؍f�^(�w�_>k��nu]R����H���,��,��'�kvE�t3c��M�y$H8����%�X��kEu"�p)�KO�20Ϙ/N�_��!?2S�����:��x��t���$Zf�"	H�.W,���+�7���v"��Nġ:8^ש���)x=A�I�j�SVQ���jUr}}5)fM�P{dK4��뽃u��<��
�v�0�*�����!�
� (��&��G|��o��CP֣�1�az�����ޞs�o�.0�l��W���-�����i2[:+3��� �`���[�0z8p�[[]z��]��D�>�=�R��Lf���D�L���\�D�04�.LSPe��9Ǖ�9ב��E�>^!�Fy��l0�D���������� �%�����V���:\S�E|Y���8=����yO���ڸ�V�>b������JE���Q�'VD���rKnjh��T|�Iv��/�+�_�>�h������±R;�o���&�h𨖈Cl�6C`B�;Y��H
������A��y|E��\Wg�1�����\i�&���=��²UZ~�үjԐo��͔�g��rfl��_����Q�G�^��l:���:�I�r���e�Y�֧Y�D�lG�YT/!���j��y����T{����jB��~����r�{t���mm\m,�b#~p��V�>6ճQ�\���x��YvvK�i/�w:q���9!ߒ��<�D|���� Zm�7%i�Jh��"(}��vtE���M"���B�pz8���� n!j�	���P�9K���ӻ���D��J0͍s�,!{�VS<4E�[<�4��R꼟7�-t��Ǽ<;g��I��.���t;V���}�9�]��:�D.5%o���$��*��H��1��/��o+����������-U��eu�@�t1��d+P��Ԓ�:���:���_���btv ��L��]��(�����Z�?w��>�Y�(W}�W9W�-&��~(n��և[2�K�B|y��E��M�$�s5{PUZ=zg9T�fQ]�۾}L���7�3��]��у��Z���G�F���u��/�hv�ƛd>���������fO����[�˅p���d��@q���$�]<�~r^�E��Rj�L��j���2:��V�����B�.��|?[�,���	�e��/�3.�A`���c�ȹʱ^&�vU���s~�7�@�FÈ[�82��X�H��n>�M�~�Ͽ:���~�uy2��ҽp��I횉�2@l�m�t5��T�`�`8W���$&6t1��p�)��D��ӏ�#_��~/V[	���rq��jI�|������_<
��z�Rv�h�����<��#>Ɏ�,����Ӿ[>lA�·�w�VG�N&[g9����-nױ�v�#�F�J�d��ri
˷�ן�M���ݮ  U�/7�Rb�()�
�u� 	�.�3�Jk�gHW�zN�^Sb�]���q��95-M or_5� H$����WY�a��2q�I�,���r�^�(/��&���bd	>~��e���ܲ柙O�I�r�)f?�w����<i���W���*�VVV�^/��ޙ؎lЗ {��\�8=޻�D����p8�I�/�I��I�*�@��yw��!�$5h�:�L�&.'m�������FQ��L7[�d�x��H6QQ��6%A&C�}ڷ&#ף�!�������n3b�I���&�d���LGp�#A���V�����oE��E&��.VcF/�r�����(��i5�C�H�E�@���:��N%� �=7�un�$��Zkb������ՙ�<A/֨j�}C���5#�> @J 
����2��=o4�@ϐIA�I!��������ՌT�L8&��C��z;�#"ñ������O�f��+[A�.P#�L��h���4����^!��n�f��!%��0�0�E@��V@��!{Qr.wA*��� ��x�:Њ)%޳&�k�ψܲѓ�^�d� �0$��&�[��sŞ��ȑا�ъ;���B>]�s	6�Y��&��G&���%Hw>��^X|k2e���=�l�"�vٌS%~��&�'ۊ��u¯[���g�ƑA+����ڡp(o� �!��lC�L�orR
�l׬f��Fs�ݤ��7 E�nϴ��D��{�Y�vj�H�J�N��"_O /���T�k"(�Y��h\��O�]h恋T��0io�3VK��ʾ�C�����%�%R>Y%���Y�=pj<��d ��2�fh�8qwP�!�Bh�ݝ(CƋ�]&���)Μ�oD�ڣ��z^��s:�tp9Q�c��}���yB������j{���і��q�p�5��_Q�eo��h����wf(�mǮ�}a1�7.%4fB�ѣ�� � \�]z��LhM�c�6
���!��Ph��x�Nt�Ǵoa�jcy+f�kʔ/#�E�n��8|'��jK)�T_�J�7 �x�a�=�^Do�t�A5�������Z��ɚhzX�k:�g�u\o�wv����,�d\\��<��v��J��31�Y��j����0䍩8�r�Sb��H��N� eW�jk�j-��i�W����H�)�=���3�,M����܆,Ε��Ҡ��#���c��mg����X�Ȇț>J_{ّV��[���!5V�z��y��1���?_O��"��2>޶e� ��nC=��mr07�S��+,��;�:g�[2ؽ��,����y0?�+��Z9�I��;7�$�~�ּss3<2\��"��OlH,���#C�e�i�E�ѣ���=��Q,�5������4���h���Q0��7��>�LW�j���R��A����g+PNTUČÚ)q{���0J?!P�Ws~�)?`���u�����H��p��M��������2sv{�K��Ô�&/�Y��]P�8��Nan�dv�Rǿ5��g���v�fł�I����~�l��c"�����;��D�j��HW��
�r�X˓��ϒ���Xp�H]ʚX����z�n&=�B[���ķ���5Q��x��h�"M�0,�ij\�'�:T��^��X�4cƀvȓ�������2�8�vbx/hq�7�`
�����x ��?B�>�zLm,C<�x!]�&'�J#���~u�ub=,��Yse����U� ��h�����ܲ�_�^�?���-�������lؓ��W��[��Ɔ��U����K��O�Wl~zx�YD)�M��$��o槊4�p�#
���w�٢b �[]����B��܄�z�BQX�����S�;ю��fp�N���ۃ:�[�2Ip�H�];�Fno�t��>m�Em�}�]���h ������n��.*��?�t���{���;3 �~T`ߜ�}f�����M:�Sgƛ{�ԆՌ���0T#��� ]��Ճ"����Rv�!�y�sg6��e����R�Q4�tJ3F�p�V��҅�#�����ߝ{���0��u���r�#���V��}f�����;n.�xD��G_6m(�����E������妯JGQ����GE�6��M[�#��>/l1v�+����v�x=���4��?�čj3�FD�����h��6�����Yן��)RO۰FoR#�X�2���X>���)p�TI|3��Y����wJ+�An����]��tP�ᕿBT#�i"���[��)�܉�rV*4��D���M����p���k����\AhkןC+�nl%!��
��͕�| !
*6�����c���A��@�1]��y,�^S ���v�>a��$��R�N���t)��!�|�;�L0(�)�Q���,�>r��f|�ws����H�j�9�ܞ�j���O��7~m-o4�B`G�?{�r�GK�<M��=�"�ލ�ӼP��i��J����-tb�O��{��gP�4�"����+��1'׽,/���-$�8���o_i{�cu���#!>�F���ߑT�Z�ݭ����~����5�U�܉�6	p7�\��%�,(���e�9az�<���{�y�R_�?�o���i�X�~SK��]�ǚH�=����_����CfvO��R��W!P`
���9�߲;
Ż�m,����7jE�&tK�FOs/gJ2��˰H܌e��'�����n���=�)B���H�XLo���
TO]O��n/��^�p���9mm�z�F�0�BJA'��=8�yb;"<�[�Ȥ0^L<D��)K���+�6ɝЉ��r"�ʸ|��ZY��Z�
��T��X��?�6:����`№���	��V	��]CʯM}u6���я]K
��g}�����W�ũ����PP��E�"��;��>*}���W"���"V�MH��s�v��st�����N��s�:�q�F����4OR������+U�?���'���lT	�wᢩ쬼�b�����FѤ��} b�#��A x�W0]�$9���?�M�����]�?�%�uڟ�}0$�¼�=�CJ|ss�z��A����ʜ�I���*6�G�4�Wh��@�,[s���(������$�<<����S��&�h��+� ��V�""��-<h��Ua�	�
��̓�Ũ�.M���RTS��儆r�w���?o@�`���z%�ۅY��wn0+ٯ�Y�I>a���m��*�)�����˿|P�:��<Z��N�	���Ǆ�g�"X]���3��4J�^tY)��f���/�����زo���t;V��	���SF�%��\ogE�Y�����Vq�V������U&v�o�����+G���+ �(�0Ƴ
{�n������/㢩���ߕa�P�
u5Yd`>;<I6q�$�%�Sa��#��Qy�0�i@ܺ�V�o�o�3��H�`EH
^������TdӚ����}a�dO�����q`K�D9����|4�^�ڡ�gF��15a������W�����̀b�Kӱ��$�����'IF]��pG9\�j"-���G�磊�Z4ˁ"^t�Ơ�����U�����"PM�"�_ ]?Y2C,��ܩ|{w3eϮ{��=֕JnY��_��i��U	(ve`� 8��C�bK�T���E5�p��іG�bJ�!ǌcPk�c��X,l@\:g�}�*���{��
�H2����Y�'9t�:���N��Yw�O���g�N�]a�S�^�C5Q"�Omi?��[��5�)�����5��&�2�Ք��u��F�CX<l�_���������[(K%1� B�W�t?+�,���֑e��.5G�T��͍��L2ǳZޅq1�J_ ��oXL�Àp�X ڼF���D׷�sz�n�
\��9���R�Z* ��FD`�͵�<�5$JNg�;w�&Ѓ+%	��>b�h� �vS|9���+	)f_�i�j��W�:�qtio�[�P��'PA�^�O�pJ��[�~���^L�����.ۣ�}�ZϪگ��g}�\�s��� 
��HV�|w1̱1h�G�c�.2� VD�V��!%�=��]�m'�	q���(L��U5�2j]���Z�a�l�"8:ʸ�l�9�uTf,�r���i@�^i�������,�;S(�=pCNA��>'�ssW;Y4�5Tױ�_�M0�C{�	j�sm�f��R�����+�,�ݹ�~4�L������G�,[.�*��/�t��r�x��,<�O/�F����}��~�������pc�'�*�+�it}bʒ�����ĩ�ڲ���d\Od��˕=���Z�m�SR�a!�/h�Ȳ��#��V'��A���ENN�I,��3��29�A1��JA��+t�E0�/�� g�|Ǘ��H�o����y��}�{S(F7#'�p���E��e@7iE`L������:�e[ww����\�{pwww$���Cpw����kν���avS��jV�Yk�H�����Џ���cA��%bh����$^=���`=諅�f�h Y�jN�Iݗ3v�P�P�ε���zt�|�]@�X1�^����[��� 9� �ܪ�A�։�&E���w��Hh��T٪FQ��3,色��˦�"���H���:�8AY��m�M7�jN��V5�5=������;�S�z>ݖ���1�g#�Y0>P���k���#�uzp�����h&�KN�eN��!�]�H���^MD�_�0=0Z�mxs�z�(���ӹ�α���?t}���������������"��{�7���z�R�񧅼{UI���4?� (�){E�c��$����^IR��N�����>ZQ= �2ꝇ���jb��~MI$�	�	�#
Xf�S��I�.���ܬ�)VkV�s�%��QG���×`�f�g���g�-���C/tX��� ���`���4�;�wC�dgH����:	�-���I<zc�v�B��
[/Q�)gs9x/4�2=E�p�7
\k���
'�2�)����Uc�7�W�-�ӳ�N��?Hj]X���|F�"E�ϛ�,M)���L��_w(N�8a&z^d�r�{���m�*�	��:E2�?r{�k�T-�0���T!#��Pu� ]��d�F�����T��[�B�Z(�(٠�N�þca�.�a��uᙳ=�K ��. +Pb��1n�z����F�?O Qo�>��>�03�1�� �*r*����`����7kw�8/�Z���3�`�Q3�*��6��(�}�H� ��8�n�x`2�h��~�K&�mixke���y�$�$�=�wM�T�F	�m��;���Li�b�'��QC�2��{@��
J�Q�}�����.�v�y-��!�4�>��T���H�]�C8 ��սI�ZT]�`\jI�O9Kwm��7 -�H��@���?t�aP7�ͅ��+�z �5�G�-c��K��㧁�����	g��	V�嵅���%�f��'�B2�9����2�&��	��R�OI3���'���+�M	;�l^я�z�(qx5�@�	U��b�_J���H����d�X�p����(䵣�%���N��8�G/�R����*����� ��p��	����:�"���/�
�?@0M6`���?F$��Ly8�"�����F)v{�_���$":��&1�����%�u=JD�4K�Ф�O���Hp)�9��b�,�K�O�+�h��o�(T0*�r��I�D�ښ��pm�X.�����H$D����Vӄ{��ޛ�8�Δ��G9\��'�� 5RN&�D� �6(􌝮�8�ge���Ҏ�x��e�������H���踭a��5�ڨ+�v�{6���6+��䏼�-��^.�B�=�$��Bh�Q��@��I4�:��_� ��Gv_� Q���I�Q��2���]���L����{���5 w�����^@��%�jf�'H�����=F��fD�hoѰ��$�`����]��Q����v�/v�%�D��k�cA�����[�"8f+5tt����y��,G�*[��_�����E���r�$mf��[AK&
�z���K �����_�,p���_�ԡ6w�������e���t$p7����"�����IBf��0�k����x�P±P◈��v��L�V�\ڈSFo�� "��A��+�޳���P��e�k�Y�d�pQP����Y}N8��c?���D�k�g"�Ҿg��0b�?�ˡ>��|8����玘��_B��w�@����Q���I�^O��D�&B(��B�i����S@��9�U�D������ �G
�C����`>��eʞj-�P�w���Y�p���G�-Z`�Q"D� �y�[i��UB�L/�)��s�-8�EZ<���j`+P�K�M�O�ڱr��Z%8�3�~4��J���Z�<@m��1��!?S�w�� ���h���9A�s[R�,�$��2�"ߦ�@�H7k$EQi�P���@�@�N?�e����- gA3�'g=\.�E�����q�B��J�Ceɰ���+5$���a�U���l�_ }ƌ-��aK��*���-�"�\�� ��@q��$�7��A��=L�5��UU����KsK�~.��o����r�>��֏TD-�(�X809�A>���,ί���Ic��	��'�e�(�.śS��U�>RU�t0�*�Sk/YF�5�N7Z7�QA7A(L%c�-��!���2~��Ử��,"$��-X�ؚER�.e�DyP���Hp!@���}��f<�����hd'f�E�y���(��@�� ��?s�B$�l �d5���<%�#��R@��y�us�2Qxb ��QS¡ x�o�z<�ʅ� �G� �/��|ߺ����Y@C b���r�!�0����zH���s��0���'�܄W�׍��x��2��9�)�+�Zb@�b-�0�wጻJ99~���1��쒯TW�Ĵ��Z*=h���~i��HH����e/�12���w~�g|�(��0��{�I;+&��rW9��!��Ӿ�����թX��*���Ӓ��/⎋:�[˦�wY�����?|�nOX:���0�Ϭr�,4r�C�� �Q~4�� ��d0�k�oc�����)�˧~+�9[�MY.�'�U�osQ�Ӫ��i�#���[>J�b~�_2\0
l�9\Cq��R��� m��@�B�:�j���:D�^F�	0Q�ѝ	 ����3Ai�C���1�:x80%�N��B#į3���
� cO�w��SW��g�DW�%���1�oԸ{4ԃ�tMCq0R�f4�	P
稰̳go-d]2��i��`Z���Zr���,PY-<��C`F2�7-@a�a`1(Y ez����E�ЏԈe�.��WS��~��]a���9!~ �H@y욅���Hc���phX՘z�x2h��%cv��b(8�ü�עZ5����T��z8���tW�#ɬ���j� ̟�<Ψ�(6�~z�ٯT��d�4���P��i2�}���B���e2�ftY ��ՀU����%��W�Z]8��A3׫����}Z����� U~}'"�!`Kw���#����p~��V��e���ܫA���|�ua7�es�a6����'�{��{���*0��5N��N�`fn��	5���!~�x_�KY�:�9Fp���S�7����2�5vZ���2�6�Q�/�#��2^�|�[��֨G����g��ң3���VjPΘ:�1�B�$_ru�OG��g��29zg�ݓXF�>>R/�!�l�fv�����A�1�Jᷕ	qƑʗ���QZ��G�-���ܖ+��=q �V��|*�Â��4��)�;Iqv��֦}��ۙ9�N��ӀQ3��^wU��Bʕ����!σ�����LU2���c�zk�u2k5�u�rz7�X��t#�+^�+v�̯F�8�x8&)��+�:lI�f<�YP�8������G>z,a�*���V���\�<*:v5���[�L*�Y�
�"����qeս<Bq���]��G�R@�4��?j��JӮ�����[`�պ���u_.��������݄�Υ~��z�����F_�)���i�.��ZǄ�����d5��{(�W�������~ZV�,sNb*�pwmBS)���$����j�L �(�s�l���5�{� G�ߪ�P���|X���K;�L�n4�� �`ΰ��#�r������q*ƨ����t���0�=qfBYҧ��(e^��?����5��Ҏ]7PΖϳ�f�����}K��.��7f���&f��1&�/�,NNNS.]0�ː�I{�����^�zJ���(�6�k�����8��_������f���fС����0��?4�II�Z�4��Gj����Qs�&})�w��M;�e�9�L Q��)h��C�{;��7���KtX-N8�B�#B��c�X���I?|� > u�Y-E��&�`I��UXh� Bֻ�R��fvY ~Cr��#�ܸ��?���C����l�$Iwԗ�I����2Fv5 ��J�cc~&�xE�|z*FN��T?�﯆�MP�J��U ��u�vDQ�]Q�|�tH��&��4φk-�5�A�l��`��#'��\S\��ΰ�'H0J�Q�Z�%�����4�P1��\i�^����BH ���_Ws5�z��y�ۯ����)c���p��\�m�	RЇ���T��������1!u��g��F�ޥ�"j����T�����S�'�1l��B�M�Ծ�j:��� �2	�xw�(��n| Q��֨�@��?
=���iO���F8�[��A�0���#����:�j��r�_<+8�vd�o�����l'&Kw4�����z�l�J��X�u�B�T�/!�����N��Q��<'���2������Y�_2��;���$�lT����_r�f����Ww�T�G/Ɣ�v�y�~��>M9���?!ޯ�s(�a�zްBlz�%������Xl�b�iii!��?*��|uȄ�~��JPJZ5��^�\�D1w������z�He28Ò��"�J^�2X��
|X�eӛ��0�>�|{�0�l܏a�FcvF��34��_2�+�&�0zPD^S��2�ڬ�N�������(	��eS�!�_k�Su�!wΰ/����C���ތ�'����p���Q?ȂG�X.�����4F�*��i@�L,�7#9
az$Ŵ�6-笱���?!�u�;b�¶Ƃ��]$rp��;p&�[�}?)�TX�r	D�R�.��mߎ0��]�Ql�u���13�*f��J ��>���0`��燶rG/h���:�Wʌ��g��r	�ނ���l��o6�$g��"�ԯT��7�=@.M�q�J��Y��؜2�SҚ��C��th�&���"�X�uoog�Cg������OvF�VC� �6_�s2 �Oۡ\a�cZ�Yů!s��+Ǐ �'7M���a":4XsCX�\LFy��������i}k-�x�(��V�S��^7׋w-L$�=ɈNԦO�f���%���4�9��ޣp�.=��4h1��ӞJk��z2���TV"�g_�-j�B���Fu�������;5w�S�2s�Hm�D-��<=�X� �B)R�٪ns$Y��7*�5�LMI�c��ڏ_z�UV��`�	����2�é�d3��R;jd$��3�`-�k�	J���0eݔ�����iHK�G��F�g���C���X�e�0�J�� L| Q=Z9���d�hy���-�y�OZo�| Ƨ���!�	�m�	��HC ;�U�$�/���vݧc��-��������4�6�b�3#7zu�2��X$�B�mЀ�N̛P.�#�[f"V?�'��	�^���h����da���� ڳ`�߾���>k�3��g%ĉ�`�dfD�B����!{Ye��=/a��:��� �h��$����KG�_�A@�o�����Sb <��&B�\�A�Sn��A�3l��GT;�+�4������+��NJ���K�̎�7��#+���}���/��w��D~b<�� ET�I��v��y�9�t-�b_��d��t�������S�f<�sm����U;W�KF�BU��fjNv�jeb$��#��-�m���� j��]�$.x��1��VSv����a6�g���>��!vх�?�0!�C"�F@w-91j��Ʊ�w���T"��+�O�1��l:Ʀ��ެ<r��K�u��L�?�41�ѦXX?
)��s�h�q�W��j4[A	h4���؀iB�`�m���t'�"���=nm۰b��������ws Yq��ڝv�l�{]/#�|�.��T~<)6�mB��ꯆ�>/̏�*]�}қ��r@?PB,�7ˈpi���֖`�AO8�������΋UͿ	���價ӵ��O�������J��v��gm�8:	���X����e��Ϛ���)""���YA��{�>a<���ySe{zC��8h����B2�N�\n�/3Y+�͕��)���;w�`/[jhM��wB~M�{f�L&Aȟ[�-+S����	��|��~j�=�M�L�9wr<l��#I�����RRZ�-j%���DVi{>��yR/�(xZ	�^��<w�U��f���f3�����e�}����
���u^<@^��XA&H$��X���B:��)��aOw��`:��"��T��{42G�����2HG[d�-���F�a��O3�E��{��#��I_�K��1�ΞΚ�\b���Ј���u@�r4��~��akv�7-�N����Ok��c1]{�&�;M����tp�P�Pc
Iq��P�nni � ���e� ��w�������n7�f�I���.MdKJ�y�h��%^ �ষ]�
V̄�72\2Nr����u���5�Q98)]�Et|E^���	��k��L�-��� �H�;�&Z���l��8��N�vb��b�d[��l|��tU���)P	�}@�89������qaC'22!`�2���Cm���º8SSNT�L<>+D�G����H�������H?A��d�^�K�� K�'�ډ�)*�ƶ����� ���X��JA�%��?������ǉ�l=�(
k����~�h���S�a7��?5<F��(��]u���],���rs�bm�M)��Q�V)�F��3��ǁ{��������E6�Y�%% �9FL��u��.rwHŧ�z��U�}��L̞Z�J��toi+��g}J:�&(K]�&�?�w��m�\��&N�wFe��-b,�a���%�ψXa�[ⴱ�Ņ�mx�eDu� sb����c�
'����WFℝN�5Isc$F�0Ϟb�Vʓ#Y��?Hy��̩��C�g�6a̴�����ƅ����֏.�;�e!
������=�	��V��	������@Iw9�9E��og��?_�UK{�3�=�n��Kϕ�����6�H���VL�Q�k��	�16N��%ciY,_�-krrrj��U"?f�2��Cz��E����M����c�{M\���rEk.)�(�;�6��mFۜ��؝īkV����e{m���&���7����?���گ)�I���]���EͦU쑜��5k8�e7$�4�Wv���?�+O�����OՖ���^ޡN
\!1�BM�����f�V��O��,R�;��6���[�Q���-:s���a*r��g@�oC�k�[�|X�#l��9Baջ�U:���V$v�-S9FU�0-s�)�]2f��6��ގx����J����<3�:i�z�����A�S��xM��p/��i��bU@o��^�Wމ��Ya�V��X>�ʒWH�o�o��a��&ٛ���d?���W����X�2'vI�9�x"ImōМh��g�r���RY�~r��W۰����,�*W��Z]%\�č���)m��>#�+�,���S\��7giT��ڵ�|W���:���
��td�}��� ��P��?�G��ƨ[dd�;���zڗd�nhN\�2��i{z���l�d֡�ݪڛ����	�k|�N�L�Cv^*ő^m2GZ��5ۡA~p�n�G���x�+=qb�̢^�)m�����u/���:l���?�Ɖ�p�p�
>i64���VJC��<�d]T��VC�k9���m���]b�*T��1�����g�e�>?CL�Z�j��[��\?���e��S��p-�(��-C61��e�~~�����3;�o�c������R)���Qn�Y�^Ah�%���n�>����N5�V��)v��\�u���ū�$�d���3L�-�@�M�Z�0)��y���+������\��o�>�0��d�L��2R����ɏn8��E����n�4��Y�4ƺ���-���=<"��γ�q1a�r��>�n�D�e���g����� WCM��)�|x;�<��M	{�^�Σ�����^}2	o�x��06��~?�#�Ll��D$��1{�Ȩ�G}}.ߏaX]�
':�ɒ��n, �y
��kS�aLW�����i�}6(=}���x��0[j���
��s^KT��G��_-�tӳ�]�N9++����}�J}�ɼf��>��f��ӆ���2��<�._q
�Rr�a[��U�`O�LR���� ^Ke�7��Ze��,��m���5���Djm?2� 	��S�ۄ�7֦��#d$��"�ԛSN����*������9�����E�x:/��؎dlu>��-3�h�S�ͰĮV7���;D�n�A|#��=��5���O���	P
:h�p����r��:EW��	�bahJ5�S�^�[`s�p��Q�=7e�п���~�oy�-[5{��/���%ԥ1s7�KÝ!.��<)����:ҫ��l��>C��|W��h7�)�֦��ǫ֚������K����'�q���V<�t�{L��}`l<o2h64ꙋ́S����W�	�e�hw#�(��Bi֛0������xɷ��R�'�v�+���N���0q�GW��Q�aSn�)H�~�oY���z�'�vk^ZSd�
����nU�ݚ1y3�S,���St�ʧ�u����j�������0f#���r[��u��3�R�DR���զg��W
	h��F�8w~߿!W�F��BJl�
x�d��+�콓I}����DM5~ I;�q8H m$���maܭ��$���5���	q�c���t�?w;7������EGV������;E�䡬�r;�_%�cs9�0����+��x_;"W��@%4�ဥaW���W��H�g��SQ?���:�[�&H��2�$��}����M8��<����A�o��5�I����בԁ�b�@��,����M8��(��������P|$�W Uσ�8^I�\���1uV)��]uP����8���T.��,,|�	GrvL��6�-K^�*��^�ط���b�X3j�E�W<�"�0٫�[��J����#��E@��MLi�u#�n�Z����ݤ"JN��l�p�q+l�<~�m�5�;)j�!��Lһ�q�s1d&�<r�����7���t�ֆ�D5�}�~�ֱvk�?r��������E�9���j���QAS;QKCEس��d*�|~���S��q\�OY�����~_�}����/�yS_s;����q�S]s���*]��x���b?I���5RZ�Se\?&��
���9�	E<���S��	�����/�/]3�v�CC6H��y���/c��8���P��.���Lξ?}�+0EI!���J��h���:W�AX�u���_�_���@/k�iVr/]@�}~��&k����*J_�/�n-[o��S��{�����@�crv�ꆫ@�x|Mk�.��e-Y��CV�B��?��c�M���nx�pR�F��|j�!��]gB����A"[���Lo	��݈������$���G�[�wˈ'�����3<)���˅�>���^���߻z��k��3�3��%�C�///�	�\�O�<]�iֿ�����Ty돜�f{4}�RZ�'�}���� r
F���0�A?�QK("m$��[�<\�xj���9CVWDBcY7�����t��&���tX�
6k�Θ.���Mqq��	�?Ze!rV��&�ݒ[��6��Vp ���� �/�m�5	Y�t[�V�@�f^�)T���V&��s���5*��q�e�V�ο`'{�ai�w>�dU�D=���O1ǯ��]��y��]��T��h	�'II#J0v b��\u����_R9��{��.f�3�������T���8�Ch9�XT~=%�g=T���覯(�|;�iR<{��LuF��H�i�����4o�9P�4G��b2�ݣQ����I:kA1F<t�M������xۍ�ɂ%9X����>dN����o��K���6n�o���7Q!F���e�;%��jH��n��U7|���8��i����ʽ:�ݑy�v>�������7�.dj��Ե̻�;�O����3--���eh�1}N��=;��^�a�/Y.T�)��뎠��m�l��Bo(!��d~�9~�Z�����]�ȫK�ѳ���W�93ȊpO���NM&Y������I�+�")|Nw�_�43&��Yοr��ê�E[�Fo�ɫ��]¢ndS-\THJ�q����W@W�^P�G�(H
��NP���d�mh��?t;bB�<��b�+��M�'m�dO|����(�[��v���;i`kt=	_�1�Wg��Ǎ��{N����5].C��	A�0�3v2z�|�RE�G�"^����8�-�2;K�d6H�O�n
N�8 ��u��p�<T�Ve�Y��ۡj�G�i7��7��D�u�ƾ9�ͅ�B�����ݧ&.Tx_E�3ًO?�)�t��IjU{cŬNfC�Ga���=t��c�
&�?��>�M)L�|��#�y���܊'xl�=���U��h}Ԇ;3ܾ��9��b����Ջ�:��w4
����9>�}�?��':o
+sqi�Ӷ5��zF,$��y����c���4n���s�}% =d�wr����G^�=/��tQ&a-{��q$�F��_l,eY�z��GZ��?Ո�pt�a�h���ū��[���#�@l���cU�^��!��o���ۅ�Ο)�k��s�O�1j�A���L�!�c'����*�h��F����V:�Dz�&"Z�`���wyH�&Pf������]��ja���Ew�!@ڪ����%�K]���} ��������4�grqL�2[%��%��0`aK�O-1�_���+�3%d�lD����g�0���3��JV���W�l�-�\\�te|oh묖�n�����Z��u_�Nk��^��s�S*��(K<��q��>gC��ՃD����)�z��c�قր��WŞ�0��j����ӱF�ه�w�%�b���q�*&�?���IG	��A��&I<��:�:�g 
��X���y)6�#�B�S�j��ɂ�f,��]�zm�G��H�Խ�9�x�Ny���{0�.5<��#R4����ȷ�6��?�|cjJȯ���o���t��[g���Z%ǅ��a�O,�KY�2��,���rX��r�?�����EZ�Jw%�YA��F�G�h�����a����@@�	f�����n��U	��O�-Z���U�3��#�v�Z�/��X���|FF�"u_��6/�i!=L�
�����xM ���R��Z6I}�	�'��i<6�if?&q!ar�� �厉̋��AY%��.e��Sm2<FؤQת�}į�)�B�j�[���a�!��5$;����ʟ��L���繆	ג������~�O�~·X�Jn��7�1�I�����8���*��H�
�`tR�a+3Į���zp}�K}z���r�z���qblb�{m��\'U�	M�ۛco�H~�q)�ť���pH�9>��W�l��7��X�I�G��^��Q�m�+1jbkzם���RB�����J%	�Z�h�:ݷr���i��t^����֔��V�����Β3CKP��1lGtz�pk
�۷�9/'�I�4P�9�+����, 9���'��~����6Tݧ�dL���=e��Z�w��k�X�F��
v��jmv����ǝ�0[��-��T0片�� J97Ci��'G{Ia`a�X�*4X����?�1r�S�^};�ۦn`��}����&#{|�1Cmw�I��z���3xߚ3��}�ϧ|L�rc�.���(�JYU��x�1�e�S"ʖ%��Y��F㞻��1S���<Izsȳr�����&`���R�#���ىt�_�����?�#��T�kIP��ΫC��zT�P�� F�(v�]Mo/�r��u��M��]���N1«�\ѹ�uO�"�+��x��^�{�9�6(�֎�Z(�����g�ؕo��l�L!L�B��ԏ�g�Ȉ�bx��I�xgB,�D��}h'ӯ{ZT �ή����Պ䋸������;B��m��W90y�<Y��y/F�Mb#���Y����[���ev�U�f/n�3��_���<�R��I�Œ�8�dE���3�/�>\�`�3��_��@���P���R���>�p��4a�sR�w�k16�X�����m�<�66����V;���v>��jz����Clo-�?v��R�d�2
U�k�αm��I�"��@�;^?��>q{��y��2'�G���$E�g��b������lw�]�����zD�6`�{pз��׿�2����*������*¼7���O��$h���TcZ=�A�^a@w]���}����m��!��R�߃��ըO���x!���ym��57�g�o��49[ֵ$,(|�>r�ކ�y4�[2҃nJ�	���˔�P��Kbi���E*ZAʄ����w���~f/O$a�K܀����w|�V6)��o�"��|v�ʔ��o��Td�n3B(@��1Em��]K����"�jqV�(���zō[��B �,ZP$�XUKy�kUeײk�}C��4fCD]��N~ǃ��맋�a�2.���| T(�y���gS��!A]�5�����F�[V�8bv5���n���8٢P��oj;9��!&Xh�<�W����<~��}�Y���H^;����1�x_-�|����S��p��5�=�q]-G,�^�˿E��+n��fV	���?��}������u��\Y��HQ#�HD�ŕ4G�Q�=Ow�z��D�P�D�Hk���lZ�D�4�6��T�m�&�%7��	(��"̊����HH��/X���rG�6�*�b~��-Tuv�����̀�����g���S�r�@i�v���G���#:�j)¤s�e��Ӆ5߫�e�1��;1b�����]�D���_ӥ��\o�vρ��F$Q��x]�g�"�)9l�	xN�=_{�gGBڌK=B��-�cڕ�cS�K0�"�H+?,�ln6\��nTg�
��,	�}�f�"fiw���׿H�P�5O���a���G����ʞF�Mwx�6��k�P�eO�x����]��dT��j2��d}p���^���?�N�y-�Uԏ�Z��f����Rd9`�.,#�Q��c �'�2�x��X�k)je���w�ns�#�q;Յ�%Fn��fSo�K���Gh!�I6��oy�K]8��^�T$9	���mI������/�x,6�SB8��s��/�@)[�ɽ['al]ձ<���SP$�sh��?܈&V��osG��K���͈KC���a-Eng���5bU��g���1#hp'������oy1�u�MaM6c���@�%jG�5v�O��%xgB�q��5)��H!�����kAj��
=��ցA���!`��mq�
[�@�cM�<���%�2N���*!-��5�Y��A�6���π�v"z����|t\ݶ���	��[����"�Ywc	��B����4���^�dg|+�6��ː5[���YqOvG�?�������OfN�|jMT֡�j}�
;�)r7.������VXM�1��_|$��̵ǓGG)�k5����~rTÉd��&�OXwW�����V�dvfK�uI���/�A#�Rp�(�z޵�,����u�� ��WI�5s_�_E���|5-�%�F�t��uU�YW���Ws��Nr;��L*8��̻-O�`���?Ҋh�~8����v�<��ţ�(�I������s[Ʒ��w�
'**�_�pG��F��X����]�K?�-��S��&����ې�8;b�\y*h�H1�z9sM�>�CExs�g�îͿF�CFF.�im���"�^���J�g���U�ȇ-m��މ���	���#���RZ�������,,�S���;�!R�XUe�BQ,ǰኘ��sB�s����ASH�H��V����J�SU{�H �:C{h�.����B7�T�1�>+�@���~̾J���K�]c�{�0=�E�ry�|��9=�fQRwHWá��P�*��^*?�=��_'T�x\;�7�<�Xto���I�>J�]o��`d3'U9����%K�)P�Fk�cҹ�ӹZ��7ۃZ�{s�!��h��~��[G��6٦��f�R}��j!]aȾKu"�Τ}"w�]o|oX���g��<d���j+P<ߏc�(��fJ2��%�Y�N}�C��^���,d_=��M�ә���$iF�3F��E�P�=�͔�{5zݟ|�wlQ�R���5�!��{��iHX�K��&ē���1��o��{��j� ��6�W�C��$�U���w�0�vu�8�d1zב=uV6Ƣ��X����%���+ۯ�iL5S�&��psJ�C���'�G��Z.V���l�~˄���x73�G̾� �$�4I��ywz*�9��lz9]1�w0wz��qK��s�I�cԳ�A��R�gce�Y%���-_�G����᪇��Eba��D�{�Y��i����DX�Ǖ�.��$�&y
7�1.�OR�ū5Ǝ�|�����B�tR�ٹ���߇����I�`=�X���[�C��6���w��T_�NM��e	V)�4L��/�mG��5�&a�>�*ms���&>��@Nw�X�I(�g
�C�@�d�L��%�RG�Zw���#Ծ���͡�Ҏ���"W�f|��$2�N��Χ�O�Jv�U#l�CWpAqvaS���V�r9K��ޭ3���5�\>�z�J2*{&]%��[���j�7;8���<h�����B��Y��h�bG�vI��{ɼp��9$�ݺ˜�;�oR5A;�ɂ7����rv;�.�Y(��3(|Rf���$u�)����ܱ��J��|���Nfa�9�x��91}H�ć{p��#/���Yw�@y~��*7�ʂ,�g-�t�����W5_��.KMs���y��m|��mr�o�M��M��b�6=��6}Y���(L�&��z���sqT-���k��av��c;W�gM�Th�p���&&p`�.���%h�J��۠QɅ~^`%ߙl����)m����_.�) d�ƕS@3~��J6;n�-N�n��WN�Ȱ�咈�~$	3��|�HN0���@9��;R
�ОE�Bѽ��׵es�$��A�O#I�I�8�i�����W�P?�Ԅr�(�6=��0+.E?�4%�A�L��ͽ�e#'?R"�#}�� �w�_adLZ7o#/�8�����Ppp�6Y���v����2��7s�!dj��Z��98����!A6"�����ڌ��ǎ���ؑI8�#��?�*Ă���+�7:��,������;՟�>�vhz	#��FJ�X��d[��քP6����Jnd�)���������v}�h��k���,2���?Ǣ�4���E���ۑ�3�n��6�2Rl5��ҍ�2����ݧѓ�(�-�m�ؓ#��.uN;9��d���˥;|���v�2��nq���ƚd�7�M�o�����m3��m����,F�b-�;��H�_]��;��4��C�����|��V��-���������)f{����NeE"�җ�{~-3�3�,����[Eg����gńM��3<faZmT�,�|�B�r�����IV�y9^9D]rH�u��.�L4J�����L�Vx1�`��MY����S�6�hu�����J��}�
�)F:(s.��u�4/��FS����K��� �D�~kz@m��R�|�-1�h����������j'q.�4�'tQT�_Q�14T<D����%Q	{�T��1~���Vs{D����4I�C�Ƀ��&�r
�yj +���N��
_�i�Ѣ��8���PK��lx3"#�S��HZ*K��X�qg+�U����aX�N8W�J�����H���=�q��7�'f:_Y��z�'�HG>��S�s�v�}��h��D��٭��m�t��FSA�1�\-O���b�J��$�
s��
�20;�޹_������##��|is`���z�I��᨟����,�v�E���݌s؟��ݖ|Hq���
ԯ[^���XE���w�7��P��fJ���J���^�(�_.�'����=w�u�w��1ٌ�JB��Y6�"�Z���H��hHB[��Ԋ���S1��B��_�C��P��t����|�~5?I�����NP	/D@D����:���tw���X|�z�}&"��]#Ƹ�Cby���������z��?7����J�<�H�k�^���_����,bH�R1�R����,F���L��.>/bnu�}L|Mo ���1d�'�A�q�����nBd>4Ǟ��S��l7��Ҝ��=�G��z?�zX��K�Ds�� ��w��(#��,�y���g2&o�z3Xm����/��=4��x"�^a��#p�+���%���>�?��1:���v&�msb۶��1�ձ�11'�m�Nfb���|�{��Zݽ�׺��:�v��>�o�iē�@�6�l�I��� ���Dz�l�΄˶����$@��+)ݸI����w�H�~e,��t	�..�-�Q��OO^��4Y
�$o�]�~�E8L������>N�CϸǏ\Ɉ��8�������In$kU�y[y����Ѝ�uY�*��_HC](�Z0��x9IQ�{�A�>0Z�7p�m�*?�@I�Қa�8�, /�O�˘�K%�Sr�=��r"��\'SU�5`L_o��68-��_)��;��4�d-� � ���^#|��n7rO�]�|g�堨
�!�a����}���`[4n��2[�D�7��1��E.ri�8�>�P�j�n$	V ��ΡO��pt��;$=Yyu�N����9���wdC91&�QP,�L��ձ��/��A�q���_�9��(q�
��6���0R�sڷ�m
6�H��/|q먑��~�1��M��x|�� >�"��*���T�!�#��7�M�29Z/�7��'>�����Z췔������h! eE�����P���g��R	�}�y�MN��~'^\]KA����������O8��NwCq2�+�ED��mPb!YM��
m�f�z�9�+�i�y_+!EL��#��H��a���|4�뉺�(����;R�ܤJ,��^��$dՍڢJ���M�*U������v�ʛ�a�f9�iv�1G<�b�H�yM�=�ϋ�AľI`^
T�	�[!n�5��x�.����C��L�8���r�	7H22q`��,o�!ܵ^�I��?�r���gE
�w_� �{�,�(I��K��&|1w2#��]煅Tq�[/��#�Q��o`]�R�Bw��$��?��@��T@n��ᗈ��S�ܰ
0e��W{��8��FE��XeZ,��\��D���X+�̤Oگ���x�&v���:;-��wlu�Շ�Z5�9��]�+�iY-
�w���|�+=G��HH�W)ƞP�~N��@"2T櫒�����a�TK5�-�w�?a5�KCA�l�r$V��-/�w��d���v�.��ө=w�JCC#�+0W��:$g`cc��jw���S���S������&���.l�ln<6ԶɅ�vP�0m*aq�zea�]��C��V9��ۃa��C����߱�����8�1�{�+�^� ����M(rW"r�3� �=H����z~I��EBc:DCr�G�\�pb���K���J�
2�m�T�7&��Ta�OdD2� ��Rʨ������P�Ԫ�9Ŷ N�φ��5hv%&�#�6��&�<TqS=�xV�
Y�R�L�0R>��K,�>0���j�řp4U�������e�{G3�.��q6�YAR8#E�U�sl�M(�5֩�| ps��� 5c���}����^�N�?[բK
��,���^4�����1�*n�Գ�Q��v�c���B'kJ5lJ����d�m�P��׆:"N7ĉur)U0��+��XLkqS��%ƶ��ʍdya���X3T�����Oa�yd�:b��l�]�\��=Y��HM)���P��ʻ���P�>�h/�u�b��K.���'E����q��Bْ5� ���&Ԗw��M���*r���Ԓ�M�_����.��ǔ0����(%Q9�IQ��h�H-��M�M���x��	�Q�p��%Q���q>�����bG���l�~�(�~�F�7��H������&�QT}�6�����Oa_܃�"L���`d��b�mx|��Kς�����R�I�A4}G7�`��G0(�U�(3Y��DY��ݣ�c�}�MuU�����VӋ�Q��O�&'������tII�_�jx�co5�3�D��Ö#Lu9D�b�)��\�N��V^�Py&�n�5�%^�����eO�.�z���KFT����"%ĶW����O��7��f@��}	��;0V��ʡ�[v��D'��{!rg_R�e��G�x�%'���X4ƎE�]��v��524�U䎎��=lrdD���ď���3D�r��-_r�V>J8���V��t#)̑�K�x&V+j���5���	��I&�H��N��5]��p�v�
�����=�q!�?�=�|��$`��s��:&R���CA��eO�,����˃��勛B5ǫ"�L�'z��K�6g�ǋ��vxPW`�{4ѱc+B<����P�He@��A-b@ZKk����;C;��]���һ�i������"����kq��}��.���(iܡ�c��?z�3�z%H�$rG>�%���^؍�bb�G��AzJ?/d�bѹ�5�U�|>���������d+gv���7H���������7#���c<��7w^z1擂p]�F�o�V�A��ԇ-HY�"�EԴ��/ ����p�׵��Qu�Un�$�N_Ҧ���](�I���WK�`{�H�:Oĺ��D�
N̂�Ȓ]�>A���|��6Iz�YeiCq��o����A0R���������+�%Ceqbic$��!�g�Z��Lw��b�oY�l6&W��S>���3x�������8�r]�T검��Duf3�6�9����<~��Mc�4�d�QQ.���R�;u��޷)X#4ߎ2��u��9�:��m�$�H�������Ɗ�'y�}���$uԚ
1��K>����eC�؃�C�9����)�l�����c�Y,ů�:�#�R6�:��	U�=�	���_��R���-��ڂ�5��ڑ�*G}��ޮF|�<�駶?5��/CA2����c�vx<�^��`��]-O���d������Jmff/"6��ng8@�e��P�1m N�p��?y̪iMy�7��Ai��Y����Y���C�l�6��=u=F�E��e��O��q�wb�*��D��#b��E���@w�i~㒐���{$!u��Jvi:v�F5������̨��$S������e����6T�I�a~ȝ���w,d[�R��1�7ng-eIp����Wi��M)E�G�FB
�������r�NOU�����Z��)�ΰ� $�ibv�ռkg��V�Y$-�o��ӊ� S�h�ܠS�U�:ڒ/��'r�/�͟�)�M'H�` Bw���p���Z���4�oGC��"	V�l��Rp?��=~����>Ea>t��q|�$�$Z��'n�~Z*��s��(�#�]�!��,�6�UTL��u�πԓL�B��k�ԹW�di/eJ���JAW�������r�9�:9��
��<(v�^�ɪ���p�YQ�P���>I�l{�_��0Upe�%n|�T'"�S�&:#�S�_b���
F�X6:���	�Y'pQ�j|�5�&���DN��'��_ƭhH�]��]?�N�s�Li���ġ[�^�VaL�Ph,]�ԧ�=�/��N)i��/n-Cl�/Ǯ�A=S�ۇ��~Z�6�RCCC������W�	I�\�Ǚ�,��h���e_VF�GW���zZ��;V#�K�zR���	��!�W�m$[�1���(X;>�)"&9��'MSM&'P�[���)�����*+\1�;�&}���P��8��
 ,C�}O��^�R�P�$w���O�[K��$�r�����B0(M��H�3�L��lb�2��n���o��7���U���?�7�~_�/Ŋ�8-�<(a\��X�QD�(���N��X\a�{�v��o���:QK��%�s�Ruϸ�/F�4�3�ɻj05Q�Oa� 45�A�%�i
_y�ʓ4�|W\h���)�]V���}��hALֱ7�6�9�)C�J�����0�`ٗ1-f�+~�V7N��>���Fɉv0e#o"��k��wI���C���R��c�q)��I��?[}��  ԮM���Q��D!������jf����+X���hv�x��3�Z������&�_$�Y�?0����/�V��Uώ��Me��
��숔���X��sr&�a��g�>ʱ)f볇����z-��QQ�ޑ��-)�Q~��s�~1f�-�`��+\K���'�8�&S=;��9ibÎ��^�FVm��A�Tl���uk,*�,�ro�o�����}cSg~����v�#�ō�MQ�_���@}5`�zé�JI^��+h��B�@����톣�	ܹ���yFXU��	-s�z��/1��o������\�v�%���zys�b�@�J���۞s��U.��;��yq�-����EN|s�X֦঺؟��6��3r ��W����>����A-�Ojg�
�d�cc�ˮ���A����~�S*E��.��좥�����Z� �� /��j���X���ր-8�9Ǥ'��m\�eB&E$�13y��L���:W�/��5����XpP�GR��*��	W塩)����>LXɊ��\��m�M���z��!N�����K�>/z�(ˤ:��zF���=<�d����"�IʌD�\�[E9����°˭,׿#�K�hp�[30�������}�P��G��m�_~C����Uyj�DKZW 0{�O�@F ɽR����!��I!b����!i��G-�/�*��T:q���5�|�q~���G�r5����Ѩ9��j���~|�b�v$�:}����.�iBv�KՍ��?vǌ�e���%a���ټR��J���Eb��P ��+��|��tﱺd#���ʤ����i� /`UwBPr��<�[��������d
���w�6e����j�$���%�1�<�������A?n8Ml���c�a��P�3����'�1���_)���Z�:����9��l�5D*S?O~U��F���Mk�AO��w؃5��DC�-���oTS�������]��W2<�i8g!���Ht�&���Vx��bFrNR��Ό��vό�|v�7���b�Y�Y�%ؔw��J56��r5Y���i)�x�%�H�僻�;QCa�l����M�w�+r)_�_L�'ŇtP%077��%�v˴���t��x��3Oi��x��1��/2�q#/Kj�^�#����헃¥��jJP�ة�������;�<�D��׏���ޑcO��������2ݢa�����'�*��ͪVU{S��R�y��<�
�����ӎ��9�4�Z�}�U��TMk��m��x$7ёy��qI۝�م��y�R��d)���bi?Z(pFwr9@��/�����������2���'|�Al堩%���U�$EJ����y��.�,5�`x�� )���X�T��q�����%��'��<I�m73>�~��cۥp���`�Ү\��n��k���Q�}d���EQK������N���{����l?or2�K�������藠����Me[��gζ��.�E��������jv��;H*�~�u�x��#WhR��/�ܹ�#XV��[��|�M�#�Q�l�}E-Y��L�j�:��&�T7W!$��A��d��c+,C��>�.z��IPC r�SYc�)1�}L����?=V�r����5��B�,�0T��K7���&��-⚠�� ���Wu�I`�r��@.��^�JySn��-��%�*�~�8���3Hϛ��(���Od`����̚*��K�K�?g^y����Q&Z��%B�ݵ/�	x>����J�����ثv]���xF|��ANf����3M�w��gd}����Q�b���a�Eka�BL ���v�v�rc`�4O�Ӎ��q���fY8����#k;A#��0��S��̯��W�y�������;#�5S�?�sX�� �*��i����� o�3=6ӽ�@��	��1O]�j���
�8RP�
�n
.}�}��N����2P�vp(���wz��
����}b��&t���\�=i()��p�,�W����&�G^~LF+ō���8������}���x�
߭�O��5���lBVV���ۀI	
�`c��V;i�MgW>]��p�uԑ���)�� ���������J��Y^���c����8��6*���k�p-���XQ�K�,���W*����zZ������+�?{U;�����/Jq�e��2'�pTO����,R�^,_��ja��G�/�'�FO;���7�3	zؽ�!�����4����[7߳���'׸U�\������B#�"$��hM�(�4M����b���&�����RǪ�� q'V��̀�,~�N���`�La�R�)'$���W�����(.���#�>�/$��*�5��;��XQo�=��S��q07aI��� I��;�5�Zv��g�d �W���\5^��Z������r��Ȉ@%nȫ��f0���~�=�gF�ȧ@�N�a����y�s_׌��� ǒ>�d�p����� �IK*Tf�9�bU�$E����*E�u�k��o�E��E<-Cr6�����wu��qpuM�\����ΖP#q�P�=�5:j�QV�m�{p*$ۏG� F�#�'�n'����j��^X tU��t� �B�й��:L�VP�-q<����1`��!H�����v�>����������Igk�߽�[?�4f�*$:Qg�8pV�j�n�;{�\�!�}����?�7�Ӿ.�^v��xE��:.Eꚁ�.�:]�ռ�u��D	�t��o
0ě�J����7����V٠�;&˟��\ɨg	F<�u��e�����"u��R_��0t�j��U|���=i~�y(G�==��GЕB���1"yhǁ'T9=�<?�t����]T�e>B���GK�p�u�c٭�� ?�H�U�9B�Kkx'$
0P��X'�{�V_A���;D[��3��U&�?��|�q��I��: U�!����`�[�iQ!��;����\}4�a+����۝��^*���
��ͦ�@(�/MCd�� �V�Ɓ���v >)i�D�8ڔX�_�d:f� �.ؔΞ�v��}�$��ǘ����˭�˖�R��(`�JJ��!]�'CC�Nwd5 �vÓtV�P������jq�����F�7]ڠC륐_��L��4T��j����ߎL�˼}�����XKv�7f���v�i�o1�f�\�z�h���c� L�Ҩ�%p��cʀ���~�\�����gf�ɼ�	��UN�����Q16y�� ��}�Δ���m���=fƴ/|dݖ%��.K
���l[Mҟ���_I�H0bM��[x��w[�J�G����)b]_h�w�/ǣb��?A{0z�(����'y�n�=ߗ�j��s���.�}@:�*�����=��!��Ϸ�OIXUUUeC�x��B��:ӑ����˛*>M���/+����W�2����_1�.�Rw>����_5tX ?��2���i�}�-W�y3uI�,q?�K�F�_k�'CaÕ��a�[�h����5�K?��¤pQ�4s�ˮ�����hvu�OOm�f�} ?'���O<��+�Y�}5|���ʇ�4ql��Q�4}��l���a�'��Gɦ�؏ ͍OD3�6ݟ��ꛛC��W�n�O�����h����k_sΏo�I�-���U�ȈL%����v����O�)��V>���z�\Mw�]�T���_ف�O�������������/������gԛ�-��ng�3�-z�-R�Ռ�G��6\x"x���%@�U<�'�!ȵ��?YoGI���dҾo�c.��VLJ<1��Vl�9���z]���?�>���5EisQ���i���f
U��Ln8�Lv4�b��W��.����Gx�\Ej�6{Ej����R_U���\bL�O�����i�wц�~a^l�����K������x58y/��3ˉe��+�Yo���tv� ������?�[jB��5
7����^Ժ�s!b6{����T��Xp?�=��4����I����ľ݇������<+�vy�x=$���s�����j��u�C��Z�'��7���`�ʦM��}�T���}烹�P��cf��-B3��!.L�J�9C����G��U���,j��zlf)g7��J%��-�zj���75'���������\T�T�|Mߔ/�r�S� (�t�-��֯޽Im5�;�����s��:'�X��\T�Cի��9i�MgB��9*��2wa[�-�NiA���������ؽy��R�B� 6��۔�ǝ%w������Ou����5���O%�kmy����[vjx�����9�ϱ67��
Fm���r焗Ox�}�Qֵ���_?ܾm x�vc�9/ƅ��4ӣa
��<������~�x���=��G��5�����q?��"6�8��[Y���j�B��$�p�8;\H��`�<�^o�gN�%յ �z��������W)gM�{��@z�h�rA巫���)j�����"^�)|Đ[���=�������,u�n;���/^i��r�`m�	�6!�\����>�Ee��D=��K���B��O~%5[�z�h�x�|켅����2ܽQ�{B.�y�V!j����i��k2�H��Hg#Ŏ�Fޟm���(W�"����K]��p@����)�x9����]��J��£.b$�t#��А���V�{��)��9A�\k�r�=e	M��M	9�'k���\������A�ikx����Zs�|�ۯP�"J�5Xf�_lqL�F�F�I��X�=�S�r7j��_F�6��⼑ɯ�
��D��o�t�WD��������8�x{u�������N��qiQ���\,:=sv��UÝve���
�*z��z�J��+����=��N>�hp�sE�V�I�07��81���zKJ�3F1}|�9�v塚-�vw������%�бT�r5?��5R���$�� �!RR�:����k��>�r$d΀ y�eJz�a���:�E���|I�!O:�C��6\�l7'H�D���1�d]n�A'� "�r}��!,ӽ������g�W�'�>"��G��E��j��M�^B�ߺV�陻˴C�#�##�7n�ߤ��WGMD�a��˻P����ф�@ER����B�=t�6�|�FG���o.R��8?�J�a����+�sj���y,�jX4���Fo�A�����& z����Z����cx���~�}���S��f��;Q,����@׵i�1��P��A근�]f����W��:��6�G�܉�h�.DR@�|��A���J��@�;nd1h�8I���VAM�����v;op��G{�F���B^�S�8��d 4�&��_ G�{�]����}�h�Ӆ��_X顁���I�1��i�8[�o����mŭ@�k6�IC���j}O�j�J�<�=s�+�DL��Mg�Bk�=����W#�T�*I�*�sZ��§R��SWגpՒ�f�
��G���3����Ğ7����J;Zf6Xy���X��%WI�^f-wi?�v�7�c�i��"����Ek�r�������*mxakJK��3����P�K4��p[)��M~��2� �#2��A|�	{���X���������o��ͦE�w��2	�N���,F�˖�#�$(�60oZ�/:x�/;���+򩗀�b9�ğ��sSO5��Nd�0���-�^�nn�\^��l�� Wv����-���c�_;r#��.l~��N_/ȇ\"��7��Lnt�t�%�~E6)_
0�0��L���%ͣQ9yw͈bbɗ�U���I�z�-�~.�:�T���~�ZL��������H���s���H}Ye�{�,5 ��E��#�}�Yя��L`g\�V�;�:9pg}������ooÃ���^8��c� ���v�XnU�4Ť�4-��:�~���	�d��y�sr�){7^#x�|�޲�Ԇ��u���Y�fϑ�&�@�\^Z�y=z]����/qT�z�[���<r��dB#�
�q�A��)����3��T�m�n��q�эq&&��a��J��7aXg���[���o���Ej6�q6E���82�<ۆ�<T�"��@:a.U�#4:i�혊�Ź����&w(���d�C�cX6xxS�T�������-9v�}�0����5����rF����t8s�������/��S�)Z��WP��^�z��|BYE���#�N;�������_9`l�̨�h��(�G�j�y"9�Ʒ�"�c�-����	�m�`4�%�5�M+ծ{� :~�G_��?kt��M���]�~t�`o2��{ 
���콍W����\IϹ4Xj��d�a 0�th�P�n��I�G������I�8LJH����4s��SXH.P�6NQY	
=���or��m�j��o�`$Ł�W��mp{Uq�������ǈ��R�?����⟐G����3���ש�`e�=D@����}��E�g�1�h?6�����a�[/�H�������[�6���i������Ծbj��^w\�m���Zn'u���/�h���F�Lt_�j�:m\%���o�eh�-�L#�� �p�(� �������1�t�������#�y�֑D;)�V�9<|��q!���K�p𳕚�Nϻ돷���a��;d�Di���蚞<%���o�ir�Ѩ^s^���<��* �O�K��� vO�Z�>�����0�NO��e��[+%�J����hHq������O�BY���!+H����p㵝f�z�q��IqR&���_A�r�{dQ?;���9�Mq���Y�Sތ�ֻ1��悐=�r��L֪E,�s���|�
�m��u��0�h�`Y�:7;�}���^6�Fx�8�J���E��/n��������6F�bس�:H��TD��B�	4�.�}Y�X:�f.h#��O�p}3Gd� �L6�s��'T��]W���S�(\;u7���T���	:�W�II����thb�L��P���e���Xo+AD�����%�ػ�(v�s��'^@d����d��Y�����9.%�r�`-Y�F�s�S9_>t��>s��pC��=�?s�[�N��X�F<��}���ct~��&��w�����֪wY�N�i(��t�"e�*�pA����^+�lM����8�w/�)_3�������]znlV|q��Ѕ !�X��Z׌���ѓ��)q�3!Jb�D���a	I�Do�GA��w�&�v=F���#M�0f� I��t5�.N�*���i��m�z�\<��.�z����+�w�ؓ���K��JZ¯ �՘�7tI��ڣO�N�>�r� -���G�v���A7�Y�ғhH�g`�����[��=l �Epwt�v hƫ�4c�u�4kT�R154E{��͋r)#� :�~bڈ;HG>P��;w򘋹&����� ��>���C����A]�H�;AE��Z���H�S�^�#�K�$�'d��"�rFF��&�|��m��锋=��tEtˤ�*�YH#	D�;S�Oy�������8S�B��	2�m�m�{����@3),JI����%>H�3Z���L�W�SC|}5���m,�����fal�������s���]�V�Bg��l=#���p�?q�P�(��7i���:|���o�+�gO��l�Fͣo2�� ��tWLۀ�(���7A��f������P=���K� /�sg�F�B�P�T�{9����~`�*��9r �/��l~J�{�׌�\?�������Q�r��VNFK�B1l��h�l���T��n���I��t�l��Bct�����`�9[(ޓ��F�����J�v:��|��B��O9m6�v]���&�^�[ x�e��ʽ��/��?�uI�3�kۂ�;?*�>���y�=�<�(
z^p[��:sQ�ŗ�Sabm�C�!+���n��߭���Qo��\=66�3b��l1��p��g�x�:�FIms�?�2b��[c@�/�Ԥ vh��O>�E�1��������ƝliVH<]n���k�[:I�r������5p�PPTʌ��`h���h�vS���G�XY���'6ʄ�|м=b���t�"��Ot��mͮoe�!���^��;;���+RR%��t�ꜛ
��+~7�J�l 2#�ߝ��N� !��W^.���7���� e�_���ψ�hF���ڼ��5���/	#)�}$��^�R��2 ���i#��I��m�{/�������F><����-6z,,�W5�*��z+�+�$@|�E	��1�}�C�-�&eJH�@>�l4�կ7[��ɴ��p�N��*y;�Y��E{%T��({�h*��o�X×�ؒa/���1�X�ր��P�'Io��gQ��4L�ŁP;�)L������w���
�����\����N����_�D+J��|�%�[�f�����	�|����@�����R�a>��0���ڈ�g����%��YM�wy�fէ�OH�#������c:���"t!Z�IdHX�`t��meR&��$^��2�U��r�V�c]?�1�� ����ɼ��%Y+dǭ��x�~lw�V$[�3UJ�Yv?��a�����7���".���A賷��h�@R����"���B�Wal+���'�G�<�������&:I̓�����B_��/u�~��?���ŭ���!�b*縮}�p"�
�){����p��'ޛ*-6����I��Ș����烅i�BӣѦ�V��\S�G���S^��HPk���,fa;���$G�Ţ��hB4���rmt��de��F�j����,m0��J�A�tt:8e���	�g���xޗ#��eV��a���^�
B$`�����݌���,�%88&����`�M�9_≾��3�T�D�c�j�NF�E́��7���}��<���k��(�w�<��Q�Jx�c�%�#դ iw6D<�D���f�'�x��K�AP�q��D*'6����$Od[ٔ�»\�S�&�k��0���ܸ��CF �n�B�ٚ����rL��W�S�ٺ@��#���>U+Vʧ[k'�[��>���;1�8�2��p�J�I�hpY5<���ր	�q�t��}����(��l�	����A��f���`�w�f5�������ώ���G��BR��V�]�����[U�U��n�������)��u\�έ�뺀(�3�bƝ}�U�d���8o:O�4��/���`�M��#�lR�Á7g�Za�0�n?�ytoH�
d �#V7���&�mk	7���C�֯�6��D_�h�v��I7_�*�R�҅�H�~F3z��^t���yu#�r��(��R r�\Ï6/�|�HB(�h;V�L�z��A�`����J�W�9���(�:�_��f =�dA�4�����fȌ���&�Ҿv�U>�:�歚ʇS3��P(�I,Ą�Y�ĩ7#�������ଦ?Z�	���B�|�hgC��M�y+��1趸ك*\�_���m��WM=��,��pv����sz]œ�F����_&\�hv�zV�Z<�o��V����9���l6]�]��!˳���z|L��R~�'�{{\�oE;�E��N����1��&(7���}��u�ƛ�	e�܈�y$��z�8� {{�?ɸ�+%�G�Э�rss�nu$���#I�@��'z�6��5��}�[X���Q�Ѐ���17����X}��c���6à>T����r��?�/X�GP%BIJ�^���I�W�j>sQ���r��Apb}�-!rJo<�\x���4o�]�XX��ܜ���� '��~�Iu�{1��c��ё#��g�J�@�u� ��J�B3g)U��>�H}ɯ����0\ɖ������,F�G�&J8W,�?6�`� ;�$���B�QvG;N�O�����f��{�i��Q�r�Btx#"FDm�V�@�@����x�`p�l��/��I�Y;���DU�ol���d���F}��q|�J3�� 0}d�\����0,�9����]H�W�y��)b?ӑ)?�)�\N�S��#.�q��x6*� �;�����	%97�?�
B�$A"����1��J?$�3��J1���e�)�G3Q�?[���ō|iC�HA�W1��͋�qM_zv,�Ud��.6�3�Z9�D�ӎ�4u� �_�y����d'E�EI%�o���f���R^O�$�f�i�:-�d1dt�D���������sg�R
�M����A���v�葔���He�TL6D(:<���	3�̺Y	qn�^��~ф�%O_g��Ll�3?�f��j��s����0�~^�t̺��^YI�g�W��h���	,��̗տ�(�އYޡ
h�uV���B��_s��Lϕ,
��Fj.F��/?��kx�Qfv��J�b�/_���� ��[�^�!�  >ߜ���� ]��C�w���}P����L�R���*F8х�Gn����T�1x"}�����R\F��K@��&J�0cR'L�

znc#����� .;� h0#��A�~ش�GaΊ��H�HsN��a���#�6F�T�W1x\���0hV�r�����>�d]���}\G;g�l�hl��Q���l�LCW9�"\%]cQ|DԳ63bY*Y�9��(X���:*U����x��{��+%��x�͝�N$�!��R�!֡��`��렞���7~�%�Z�od�&�4ZvoG�D,v��C8߯cX�Y#�u[ף ~a����%��q�.O!�m踉�n�`��߂ �-�u�G�L�s����j�s�j�w7��G�� �>�&X8z:L$`Õ�Cz0X8� '�z�5w�l�N���x�X���������h����V�3:߱��ɘ��:�R	�"�����h�m����J#]I�RiƢ.�����;��UO(�#ژ�l6��Iǖ^�0pt��)X�4��p�p��BEΈ�n�y�nŜ)&�&��e9��RX�/~��$�Cft�p5䋅�����?ʉfS�Kn��>z12��Ն��;�D8K\�ۃ f����l^c���HJ?Rl�Й��BG(`s���Y|��l*dn�:v�M�qh2Y���5_��51۫�	ZƂ,�C	1���מ
�G�r����Zt!蒁p�^>U����n� A\�����"9�v�'1����Wa����
�0G�!���|��������hX߁�ҕ�'�y��x;E:�jN�""p��֟�W����2��X�H7h����Z��ב�m�X1��~�f�D��{w��1�<�=�)�E�͞�b[�������O�4��������zMF�z�ďBD�,Q�1M�J������X�b)a�2]
��m-������'1�l��>#v�$955Ghw����b�������Q?�,D?A���s��=1y+1l����4|�H\��|t�%	�a I)b40�����QG��د��7(;2J
�*v��AW�F���f᰺KD�Fx1`&.���
�}����G��@#�P� ��?k����P��e`7q.�;1:WȢ|�$@BY�o�n�rz7����_�.l�N��s�V����o�4)&zd��Q%�F�!����#V��.���KcAr� �2��E�@B�p�i�e�����1q���Pb�Cx�_ y��s�(B�u����-����������Y�#�]������s/X��s�'�!�����}4Bg�(�m�K�w��A�QX�!da�A����W���,�`���|(����$A1@��K@Z� 0�~�%y6�`�
	���̰M4Cq�W�������əq}��H!�Kl>@�kQ��^�d��N�W��_s-�ip=�w[�ߍǂ�WX.�;!Ѕ�5Y�����2$�Jĭ��s�p�q3�GO6�1�~Z���n��f��j�iCk�	���uo�(��Ӎ�5��Ɓm�K_�g�8PC�-�iݺ�hK`7]�:�Bj��P'�#y7�рg�Ǝ�X˵��1�(,,�tp'�w� m�0��p��������i�"(�d0_"�L����	����3䯁�R�ig
�t��>�֊mV�i?Th X=$��PE�J�|5��k0#�<�T��4_�璜) ��|����a�6±t���1���D3'���u.�@����2<r�kX�_����@2*��ۘ�ϻG��F!��^<fpQdF���{�f7�<8S{�{f����g'6�	����^�bz�n�x�3�Sy NV̞G�`ɴ�z����ӡ6N����Uמâ��t몣��@�N;�aZ����l�O�~�Ue;�����P���
��V.V+���$��U�ʚ��Bz����r���fr����pWm�<��U#}!�I;�.mR���H�=]cc���4dH!�@��hH�,�g�9K�:m�=G�=Gg�#<���+Gp��3`�q���w(�*�%{eq��(��	˴3J_���P������n�[Z��ϗT��+�[w%���g���W�p���g
F��x�f����J&�C���E%i�յ�XZ��&�Pdt-n��x���N�	��z�l\���I�`d�YW�fԬ)��	���R�)n��ݵ�ww���.ŝR��]o�ݹ�wf2��sf�={��}��$�0��ǎ��B�Q�3.�9\Yxi!����Me6���/�sW�!�[����� /�6`��(<Vo������ӵ�"N�g#��O/eg�?k��M�@���BX�nPbê�Or �I\q�f����ONM�r���=����Y�����x;SB'D��i�$G���H���8�T����qc�I�1;KȓRL��۰�mX�S�8����+�+�[�Z��Yʝ����8��v+{�	�/	w�Y�PW��#���W]�W���Z��B�5~<<5���hp�2E��\J:�N6H�_�\N���q�\t����_��NOK��a����=ƔCb��?���p�q1�|D��_�~�;.\^� �{ݥd߸��ݶn>k�	ֆ:�$�`L,0�����*h��f���6�?�lL����Tԥ�@>��N)�@��:�!{����ˆ��v�z��AkV��$i�H�&���WU�WW�' c��D��w}.{�!�?��`A`�a����K[����=�+o4�T�_���%�B�����Ϊ#�+��v�8�٨kl���_wn�4�i$#$~����;��y�zܦ�h/'�����]���ёY�2	���d�v~����"�h�i��i����B��A�R5:8�e֢�g����q�g���tF��^r�*Tb"vRd9��,�UT)��<	��wO�hg�_�������׈㠽=�P��a�)$�Q���� �#�d*��XT����ͳs�cحu��5�����j�g�?B���߬����6���N�A��I�4�a
z9P� Ke��n��@���"A?�PF�C�A�W�X�}֫��K�|� �K}��(�H�/��� ��f��;,AO
;Հq3�	��3q\��:d�=�[��Sٴ��B�n�"T�c�̚�����o����[�|uv׌YJ��F�z(6ꈞoĴ����}`��u��\!�[��Ӟdj��.�mWG���	2q���k�QC�B�Ob������}��I����=�l1���H�����^�B���㕷C'�:u�[x�@%�%��\w�X�����֋FҪ*���0�)����ރ�����2�9�-�,�+�R����!C��iBU��#���ZײB�!ż ���т��.���M�{�`�ݏS���%�sy<<LnTX�6�H�6�{B��W����}_0�=1|[�G����#��u��h��TP�{w��ςa���������Pc��DGMa�A��"�ڱ�	I{����n[D��ۚ,��ֱHh$0���OkǞ�9̂l���� �����k	������J	��yNui�Wyv�7OI:iz��X�K+�,K�S�nSr]��P�@�46�QOҚ���/^��j�%K�2,��IR�h���,'.�U��|=�M��H<�H��������oӓ��=��5�������Ep�pc}��8H�j��B��g���7��(���ߒ]k=�������׽ɋ�]f�ay�'�<�J�?�e�e����E������JP�V�_�͞㓣DRP4C�H����t9E�L�~�6�2��\�+���A������$�g\�!��*�gP ѷ��_�8\��|�h�Jh9( �\�];iF�!XA��5�_�����oj)�6���=��U$�Y)Z���2�p�ԎD�
DS/2�F�4fd��#h�^R��Ľ��hV��^Pxl�O�I �4Kכ&	_�0�&1��z��HE��@�Y���B�*��,f�O.	� ���#ҽ�@�	�Ɉ#J-C�M�w
���&~э�D�Cv!�R��W���`}�x( �c�1�R'ʨpt��	��Q ����ٖ�I�N����l8�G 6��i&�h�R�(D1h]T>O����܃8�p)~����_PoO<"za��U@\~�-,(�G���������� R��Nb�3Xnz�>j�+f�`��p�;�M �*l��o�я���ظZhHf/ql��(Y�����{�Nj�<���^cqT� ��`�QP�ke�%���q�������wl&C(�����7��Ǩ��d�4s:��ȟ�4P~�1+�nfP`�B�6�,����и��,��������C�ڀ��b���s�Z��.�����*%°Tk�<��Q4�����t���ף�n��� �?I�-۞� -���;=U_�z�~�>j8ɟ�+K.a���*�@PǷ�az�׎�2{�`?J���|c��p��
`b0n*���og�I(1����|6U;@��Bp�����	�c_7L�i�Z�� w7�C/��P���[�٪���-���X�z
��v�����s8��������"=�|���8M<�`Z,���)�ߢ��q��C���S�&���i�>x�seƳ�#��%�Zd��E��^�|���W�}K�Q�/��x�R���E����_l<Wg
׋��a���8(���eab���� ��v���˧�YB����x��B(�p���^m��NX����s�B�`+�x�ӱ�V9��.&O,S0R2C#�;Q��"s3J�����|��_��(��HA�5j#�&�� C��9�L��(�T��=?�3"���Y ���	FVivp�����jցzGP»�G��Y[5��$B]u5^
�,X��h�.��	��ѯF��#�AX|H��m-�� 7i�N�LC�d{�a2J��!�c��|�H#k[�2Loo��M��lr&��qcɹ�rKo�^�Lj0 �^�Q"i��`�	8�ɽ�d�*����;
�]%{[�XZ+2���$���?Y��&�7m����#b������Z+_"Z#��ș�'_''�I�W;^7�7bW�IE�g(R�U�N�@k�2��7觓�P
�U��tZ���o��
 ٓ�c���-�aي�/�O��_*�h�.����j��2�ˉl��s�˚եɷ<n�VJ�~�	�jS��N�Ř�IH���s�*z�D�C_���6���'#{~�3�q��r
0�R�L�r�Y��bg�t��g�v��Y��Q�8w�ꅓ�th��.R�@���yG�#:�;l�e]U����۞Las�0�r�w5z#�
X����Y�<�<�Hk�^EMy�9DQ0@����,�W\
�\�1_x�+e�E"�@ރ2C�����j�N�n.�(}�r����Q�ͩ���?�=��v����1�v�Jl��-�����e��U��1r�+d�S&���
�5}�2�D�e�&9�r�@Ra��:	NIp�� �||�u2���Ɂ����S�D%`S-j�a�gͧe�O�E�Fx�EAɧ�;r��V��I�EW���C1OA4V��f8��'���{$d�����'#�� ��	J�X�1���;D��]~��� ,PWq���.z>$�<?�!�-q�T�{�t�����S0d�&���U���t�'�(�.w�7OB�����b�eu���97u�����d*d��\���Z�Q��
�����'�e��wZ2�;ur^CO�ts�z���m=�_n�6�W����|_
�j**����k�/pB6/��.##�U�Զ�aܷ�=7��T� �t�恔�<�vcZ�=�:���x:�F��	���hNb����?d|X҅�I/D��R�D�d7z���{{F�W�CY�����:Z�pŭ�/��F�����w�╲ZPJ1��_���$�C�&s��vBL��k+�wwR��Z!��vT�W�46�ų��&���҃��)������!}\\�. 6�Y��{x�Hxd+,�wQ.�!��̂@L�� �+�N�<��p?� (�|��ed�ut�0�Fꗫ�e�8������\��{1y#�U/��Q}��)
����>��8����"� >��I�!�_uűp�`⒣;�G[��k�I'
c�ɐ���y0M,�e�K|P���H8�=�(�ÉIwr(|�<�����hj�����V�x-�w^�ՀF���|W n+s�j|a�iS�R$���-2a���3C���\�'��)�z�&�T�G����4J���P�yhݐA�s��!~:�,?�q��sgu�0������K?���@��V��=M��Fh��������\?�����y�"���U,�7��y+[^<Y�2E��
ӿ]m[�W���)�"�B�I�@��w�#rޚ���,@��7i����R�1Oᵥ՘b^Qmq
���o�� ;W��HdL��9Y�A҈�OA~�S=��
&�d=E%c�B_��*��Ά��C��-5@�j`l�����]��E״l��8�Ʋ�S�_1W3]�2EǨ.�{����q�	��>�o���8WJ���b�zmn�K��4brol2T"���V�m9�����:�d�_pC}��%�bn��QԊb�NP���G0OE
�-�n���t���M�[.!��5�;�w|++����i����\Kꏶkg��!���|m�Jwf�	$U��u���b��đN��a����uԾ��� �[�˪� y3�T-/
�@.s�ct��=1��"�����UF�)�%���XU�xàF*F��!�fk���}� 2~������d�bM}����^o�T`��F��OK5���KV��ws�E�Y�� �q�k�*�F�!����<���Z�$�Y��F��|)��s�.�`���MPϤ���'UM ���z��G:P%��\X��Gu�[
���g�G71nz�ȼ�f�a��v�+�h�t���3a��[�W,)�0>Ǣi��<�։"w��������/�1�h��cM7���y������Cw^�>�i�V�
W|999��v.TzĶ��c1�{�˸����{����.��V�j~4�/�q�"+�*�/yR;ë�*
���+�	�Z%��@�v6r�AO�bY��sd,�J����;��\��&J�e,p�=|���m-V����Ch\V�ng�h��;����n�E\t�Ek(�P��i�t/���M�`��D$'����������%�U�n��y�Z(�ޔ�{_ᬩ%�ԏ�72�My��p>d�p�ćƇ�'�����'�[�/��a�eQ���IƧ�m�`g�G����R1��[�D���.�D{k����~P�f��Y��7�cN}�/��Z�'ԭƛ嶽/�a�1~S��HI�_�2-dw,ա�FY��kXMei,X�ۉP<wg6��L(��J�bN#$*ᨻ.")�]�撵:��Vq� ��l����!���U�4G�f�=�y,�jX����[M6�P�Q;](������釉�!�c�f�PM,,4Qq�*�c�����{w#_tl�8�$.������0�'R`G0^�5��Ol�_�����QQ[9�ZS��׆��^:z�A�2ZF�ON��1U8�b��[ּռ�>����!�IB?�;k�d���$�����0�j5�A�m������ӓ���Z|� �6
𞱛3���Ӵ�\O�n6ď �/�hV!�6m �;�z@{*F#΀�:HeR
�[׎�R��4� 1�qB��`��_��������|�[�i�:���z�-`�_//��b�1zO ���� y}�G�~��k@j�J��.�6om=qC�	,x��
�A(�^��]�O����3�,����V�߲�2�2͝�v��|c�]�:9��<�%s�ب��u��Z�{z�v~��֜l�g���/���@�V��ְE)S	F1d-�p.A(�0�(�mH�w��D���/�p)�E��;�B����`lL"l��j��yF�֜Zu�PN0nx�8Mc'��k�)J�'�Rm$�x��%�-��i��]e�M�ڼ`A�2�F�`���n,!m�W��0Zo��ǧD}�7��I�j������#�6����KzbINV�0t�����x}�`u��t�KC���Xc�p�	���D��D�U�_�k��u�+6c o��bY�"�%�}�j�h5���]���Ť�˨\������G�9HlڟɔK۳RC��5S;G�R����b�L=�V��{>������j�;��iC�Ť�=�ؼ����Xv-�jT�w!�����xj�/UZ)�7X#A�����M���`��u����B����oP�l:{�w~D���*��j.�g�R����{����(���Fb�z��c��W�SIU��ߡcR��BM�z�ƻ�mD\�&g6��n�)!ެn��H$TQ? cR��x�AWI''�r�@�p��*�B��������2�������l��&
kk_�B/:H�Ck�h����F�P�:�R�@������ls>I� �m���q�~P����A=[^V����Π��g����C�@�{W��P�t��Tԙ�$����V���L�LDK4(ϐ��RP�k3L��-:JTa7�WR�o�e]��Գ���H�&riď�4i=��ʹr������KDQ��"�v̭�ѣ��T����@��*bdz����#q4�z�����
�9Y4A�/���`/
T�c3�X�s�n�x��w�nH����AM���|�}�/�5}y���kk>��-~,A�@"���%���h�-ΈR�-�u�p+�h؝��n��MItP�.��!����F)i�A��B�4�4�Ҹ��"IK��/
dH�U{1��*�O�kL�({�$7�(������NNX�Ny�W�>j&�Q�op��k��PX�*��O�=�P�i&�,��gm|$e�L�͖D4F^�9o���u@�a
��:�]�ʾ
���-��9p.ܣ@�1�C㩊l���H�sU/[xĢ�ݗ��A<O�Ε2Y�#�w��3AF�$�?2pT��!��1�g�`�o~��t�W������щ�õ��iO�1u�{	��_6�r�G�#��V�dpFzjϪAͱ����C�і��RF@���.pF�6��,�"���4�'6l$�7)� ��Mmz�4��!����q���:ȟ�F�:�s�`8v�l=�nI}ϧ.OqY�|�J`-WI�2�;����(��E{�lpV?v�ߑd1�`[��̮fnI���ܦ��]t�s0�TI)����Vۯ�����M:D���Gq�{�~�p<C�W�$�s|#1�Z)���9�'L��
�C/I��/zI�
��*??�5�c��'�7��XQ��mXY�C��>
S�R^����Q����<�
�ջUX�j�P�k�IJ}��.��|�Y���WHY��)��� ����vqn�Q ��"�^^,/��J��Eʼ����p&[�,��8*d&]��Ȥv@M��������Q� ����-�HPD�fH�n��	g�$�Z�0vk������ jp�@�bFSRc�E��o����,c��wͷ+�Z���v�5AF:#���4@u����L�2�ܫR����.W΅���{�Ri�N��`��1F I��=�[G`�O�pT�1�*9FX�S���َ)�/[�Ѻ+W�2�4��&���;
RA7�<Ak$�R�Xð]Y�*Xp�x��'�$�wB�X��vx:��0ξ��0\�1	|����i㑬>j����dϷ������@)c�E���)�ާ�\�)F�a��[[К/�0N�A��X��0�!��7?���T��~���
nI�H���$��KL�Pc�����e	����;�"/�UI]e��l�7�����Y�>��䉮a�K�̑�ǵ��WPݩ+I���05�]У���փh@q+y����S|7(���U����v� �/%�<�5*���Oܦ��Z�!�^���[}!��y��p�{Ә\�|�dh|POp�$.��;Wu5�&H�0|RP�i���8��G���.T�};�r=E#.��1�� ����-��v�$�Y����ڵ��r�֯��2�����-~j ��Y{��||^��!b*N#�������/��u�o���PÒ��O�&GEU��]p��D��Ll�BF�M`+s�����kZ^��z����� �Rq�_��ҫl��6�����cqWή��+2���K��?I^�.���h��+I�,�1�]<�兑��G6�;��q_�i���`��nCdv�:r�,���n��3G��8}ȩ�����!i���#����!E��%�c�W������<L�&�u�f"���5�I�:ݙ;@��щz�T��w�gD� دִ�ҋ-�7_u��(c�vXh-ķ�tX���Z��;�,M6S���#h�rldcz{]K����1��.�?"�y���y�]�e�QWW��&
�����D�&0�Kc:�Cq�����8�#��l�E���L!�����֖|�'�=�-o|��)�:=�y�]9P1��O�m�$���)嗃<�p��q�f�|�ʐWSY'?�������uy��	�_�1��=B��b=�Rzf^c�y��{� h}^I��,O;o�S,[�2c�ԗ
��E�L�n��OP�^�Kͮ�m�@��/��G[���B��9^��w�E�ٲf��{�7|�H:ko��ml3�������5�� ��g/S�tc��XЀ)���v�^O-~Qj ��C>��_�8�X�i=E����V�G�$�\�L_�C$�	�V0,���*�s�Q,�H_�O6�{���>,04,s���H%�\˃B�*�Q�����&��[��}� _��X�A�X���b��[�cn�{�%$���N�iDa�]��/�� ��H���$�z�A���M
5��8?��q?w]��>���b���t���G�:���0-�*,A�(*ؼ����:��������P������(2���n!�)�9���B�w�y���8�����*a�?z�N���1�W�[4hl���-T�nv��;�4�Fvߠ`hE�����jɨ�ŵ�!Q�W�i�A�Cf-ٓ�ks�d�
�-vm�hz��hX=`��t2�XO��jZ����bIO�j�\�9�ß(��׌�j��z�V����`�����@k+�qĶ��Qط�ٯ��:�����ġ��*�ۚn�M���h�:���3�KD�*?�n/�-w_`��w�2m�?tǐgXQ>Wu��#��;x�p�=��P���1��&�^
���4.�tSw�~pjT����=k�����̱їr�jkwR�Op�	�'V�.�= ֯�lVzq��>�Ō[�Lԙev6�J���,�2�8���E�V�]<�������0��n[�ZEM�
$}v7��E���<A�F���
W�0A�
��u�9\?�V��#t�A�"�/Z�M��R�w]�����ҵ��j����F�q.�IK��M�"�yI��P��\�Je,������ĥ������"��gRg����VT�q�
��%k�ʃp��j?,�[F���_4�~�k~�Jq^柝)ണ�o�(�͍lլ�̈́�Vb�3�'_�<wB;��?7	�4tڥgt�}��W3b�,n�@��W��M�ӽ��
sOw��lw\���p�F�����&��#�K-ʊHA��C���_��\1�z|��l��y�өu��3K~���L�x�F�\���Q�c
�Mo�?�!���?r�������D�UN�,G����l'���&���UE����f���9=r���S��8��@�\uXW����4��I�z,�_{C���� )�6�9��~�{��u��E�ɩa��Z}�x���q�{`�U��_�o��]-#e?�gٸfc�r��lR�&0�&�kK<��D����Ue�������>���`�Xq9� g]��m}hvl-rv�s�fY�1��J��NVP�6V�E �����cȹ-��a�[����й%أ���o;�L���\�-�̧
�'���/^~UK��6�δu��[��ut�J�0���)/�ߊ<���_�ߎRNJ�K�;�"��T���+�T
"�ϳ�j����v7��4����ppI�`B��^n��ƜTc�L�2N��=���zt7�I��b?�~$oz����Is��5��j/���C(���s�[!+ӳ�vn�vq�ge".M���K�F�k�뫃H��"� V�78ӏ�B=cH�P2u��Ƚ��$�{6�0���t���g"�k���u�'=k�Iv�Q o{�PH�#�F��QCL����$�W�op>-�]�"�+���o�d���f9Hx����{T����#�ϙSlG��t�^���O�����#"�z�/3Qe�b����oc�.�A55�Y��m�p�aC�.s�	���/�0ȑM���a�dc���H���Q�6�9�I� U�,q'�=ܟ�����4* $k�#�e�eE:�d��S�Z��V��\�X"Fv�}�.���}`�$���PT*�F����5y&�MR�B�F�l�t�w�e><��kk�ɕ�
���G��9>�$��J����tc�p�����(�YH~�L�Y�#��8\t��T�l�J���r#����ISNO0�@xd,�R>��^�5���8U�����Ec�*�R�S�f9r6����;���Ь}�(���^��	l�nO��37U�w��;�imf=}�\�~Q3�����j���c��qx5�q*�E&@�Ħ���^�ZRD;����&G]1��~<}�N<�Y^�q��S�,uFVX�� )|�����?ɓ�B������+T��!�w 
�[3�u�|t�=&�vz�8k5w��d���N��e�,�|�ߵg^U���n/�U?�jb�뇂ܘ�Z���cM!�M�B�]����o�×>��f9�θ)��������[�ވ�|���
�M���3����V�r�����&��P!���֘k�X���ŪI	�Dl�E2��)�@eA����=!������<��lqu��۱a���mo��]��%��ț�&��c�D�K
��/������7S�4\�a���TUK��3�yF�[w����3�䨂���Y;��3�Q�ޗB�-��_��������گ-����գ��ڵT
��W�����>3!��6���bX�v �可�>�Č�H���
^;#���>������
�	~m2���2r{:<��q�t�������I�͝��T�-I�z֜�M�w, �Μ��Ϙ�CC<�m:w�A`�ʆ�
n73�]3D�,޲������܂� �x��e������z6�b�'�n�[��pQ�լ�غ�0$��&���@���&�G��T����f��<�i�Z}$��C�����G���p��)�������\o�G��|gE�I���ٍ�n�Q�+6Sk����u9l��R�O���]$d-^Y�K����ͬ�%���X����2~L�\��Y�љ1��r҅��+[+�(�t]��(���c�b��I����Ñ9���c칢J5�sh�����U��ߛ��v��c8ǝ���%<�Htجmj�\�͌k����el�g�C6�u�M�SL�I��>�D ���:ڧۚ���T��zZ(��U9Y"gY������s�����5V%i��� �::�d&M}0b��?<�ɧ�(�?�z�%�t[I� ��\�kKC�G�5�ȏ�/2�z\d��ߐ���y��)d�\��F�Ӣ�,�_�l�C��j����|�͍=�����JV6^��Ca`t�O}���{���lw��T�]�	����~�!�+3�	?~4����l��?�ϻg6v��V�7��'���Z#���w�l�����X仨mk�w)ň1�P��]�}4=�A!�}M���.t�[�Tz7=�dE�ҪT�J�=�9���s�.&Ʒ���}
\۸�1��Q��k� Y#�ؽ�_�裎���}fl���Z[F{p`���Eյr��e�VG?�2���N|.m��6,�t�c�{��G-͊��	� Zը�\��o~�* ;:0=�w]W[/�ZL�k��mFc��L��4Ҭx5~�L�x��C
�H�z�&<ї��g�'˾��H]�R#���-Mx˳<eE� �hVcp����+]�E;�q�WQ� �4?[�k3�jGE��F�J��������61L���뒹|w	_�L��� �~~�f��.q�,�6)����y��U��;��/?�*NNa^4�{{mY�t�1����?z �f��I};ܩ5�,���'�>��P�1۲�[��4U���8����.Fܿ�	/vbs��r셺(�?�;b���e����2�JI��Y�7|v��rd�
�l|�����5���>1�o�ˍ��E�J��$�>��6���\��Ho�r@c�:�/�j��Jꈿ0�%ᤱ|j%�g���kd�f	.y��g�9сM���S4���z�-ET���5�gl4
גc�Ӄ��S�$�P��#�~�9��a�<\�1�]e�Q©�v�E^!P	Y��E��z�������q<�DAz��z7A��jWhf��D q�{�~@uI!0+��{����%�>R�ț�N~!X��4$���}'&�|���|a�l1��*19�ě�B����A׫s���y�����r�'�;>	|���}�?n���O��7��;�o�ۗK�Ң��*�E��HP^��F����ɪyy�R�T�1���c�W��&���Yw����0.~g:�J��Ȓ2�� ���ٝ�_Lp�o�J������]/�����v^,y�Υ������;q�}]]������x-�A,b���>��W�j�1�%�����j�=-9Ҭ�Nr�8�_ 
l���]o�:$p����`�{$��a�y�U����%�y��-y9�H�6-3t�Ùme��v�WEХɴ�$�$���1Jy^ۆ	��3	y��4��=�ΣN�Z�\L@g����r�����&9���ޗw�c;ĳ?���s�58�qg�D��LXL:�^���U�g�;/t�E��
��Ҿ���u��? �ű��Q{��Kպ@pZ�$8��g��0���rv~�-%�T6_"Gs� ��w�����h��T7��x;AV���A���]�cnEhP�ag��Rx�kj
25� C�ŭ�a^�Ԅ(�G�iz���IF����� �B��;!~�8�_p2��
�i#+��k�����8v��K�B[�VB2!��8�<+MGq�.t��d���^���~�ۚR������YkSvwͩ��ļ�-a��r�o<_&�^l�d�g��g;�2�����`}^�o�V�P�M�߰��'F��a�/FO�^�"�� V5��� ��''G6�Pרn�W�����
�������c����k��ۋ��󳳉�wZLۋ}(��O�u��;xR1�24�k,��Z��a��x3�k��@gVw_�{W�fa�̤�n���/�j�;�ۋ#Y����#x��s ~��v�4��q�v
_��x��������!|&nͺ  ^�P�M���ݛ5ş���ӈ0g��] '�>7�O��Ŗ��
�����ˀ��n'WAA����Ɋ���*�(!��Ѯ���{!b��""!Sq��w����s�c�i��zǗ�_�Fn�]D���*dء�0oI�>f)6�ǵ���X�,F_���,fFSb�.̋K�pJq7�J��Ϝ��V�4/6�%o~�_� �DU�z���T�q�\����T��<��M�ڍ{%�o�ͣɧ�q@̠���,
C���dJ�Rd0ۛnyD>:玷۝fX;�r��]�df�r(�I�u��i]�x��\I���;}<wՊ0<���T������D�s��;�-q�F�D��T�c�a�]��0�=�g�1�3�׵.����o���~p��ꞣs���b�Oh��o,/g�5��\=]���ȺF�k�)m�5;.�CmȽ�M��>r�����(��p�2(;xۣ������������I|��S�����*��w�s��������0nsu���G��9I�=5�2�"F�������8�<U=y��"�alϜ1ꥡw;فW�NG���sW����78�)�����e�O1�E\��0�Ow�P_=���r�\n�7��t,��%�[�L��ت[%�L�R��ꓫX�gt�_�{X���v�B� ti˶�� ����)������_�}{�|�:�N�B�GXˆ�*����́<԰�mG�yć�4�0�������@#��۝���Z�
���Q����m�YO��sdց��)�� ��n'.�3� ��Ԑ/�C'�1�7�՘�Xu��$~12
2�:��Y��x8ބ���b����L?�;'D���Fc����:7�K�U��k ��r��Y�e��(�����X�uP'���6ɏ��^Pr�g��B���[�
;E�B����0d`s4ib���k,E�{<ק��̍H���=����N�y�w�d���=�K��L\��y��k`���4v��+�ݚ&��u���R�&=Z""	�A��d�i�7f�(�<a��'�sݤ9�4�%��hH��nQB玸xW�;nQ�x�"���,�����h������Q��/˼x]%f	:�����3������^F�p��9;����:�B5:��*�/���/�������m�4�(���g��J6�e��S��=d�{z=U�����f��P�/K�v^w����� ����/^ʄv�����z�?���	�� ����#_-���>�m��o���\�X�m>7[����dG�w�ǂJ�~WS�b�'V�nG��8ěj��&D�y.�����u2��pt6l�]�����
<Հ���.�+���O����8�n%��4���QO��ݑ�氟rS��.\���w1�D��M�*�l+b�s�����i|����R*��H�j�?�ð�N�I~W`}�Z�gѦ����4���z�8A@��O�ű��K������i�Ѵ��C�I׀2R���O~�[�M?��������b��
X���N�%|sMy�( r������:e:�<,R��]�b�9�5)!�O!J�oõ�;�����4������lҜ%K	�XQ���IR|�a�
, ]��R-Y_ߊӖ>5�s4������j)�ɍB��[[M�_yJB���`r���x���1|嚓��䴞Ĳ���)gl�����F)�aȍ�7�AV�B\)A����rT�wy�o�a�@7<�3c��9�|�x���vO�FWjދ�օ��"���@�JVB$WB~t�	��ӛ�(������1���
a[7XSC�I�
��=2�{�ã��1��5e(6e����z�ΔVڷۊ`�eV?��Ʈxi�����`��3:����́L$��߆-`�O��S?2A���	��t������[
�=c3Y�<o˛�?ڸZp}�/���Y8o*'��rb-tѼ�W%؎��#��=l��*��p)����zm׼?��hE�3�y�O��7
�&r`��?܀<Ə5�1M�o���{ͳ&'���O��ԝ ����u7r���H�gb�v�6�����`�bo`lBBD�Q�;{��)Nc���D0!*'�Y���H:WHSŊtu}SP���x�'�(ķ��=��� o��G)GD^~Na���AL%T�ghӇC�w�8E���)��ה�u<�N#�< ^�0����_@%u�jM�c2OP�2�w���]�D����s�������W~������8�f����w�c�?��S���M��Zq��*xi��u&ʑ��Y_���4��z(I컃ߦEd�����Gx`+��ta
E�ۚ���m���o2��eĐn�����E,�7�i��8ׁ$���_s}1��T��e�1Y��o�$nR�B9���{"�7�\�bY����ⷒ��O:�؏�"�Ej�N�)I��������d�H���XL��H*��l���}� *1/���pA��9���Y��/�]Z��aY��x���=ʃ@�,��Ҏ�mFRRVj�R����`S��|�I=��"�\`=ڶ��L(�<����D�]"�
g�$��<6�ʻ���]�ɢ֠
���t��q���=�����A�(���<eAj*M������U����y4K��H�fۏ���v��B;�؉���f��^����;<T�%��0ā��Ōm�����T�����J�q����}���R��t#V��HK������NT~v�VE�8�m`0å�Ц<�>WS)'���KT�@Iv�P�b�G��M�*.qFR���/�qM�����bi��ӟ2"k�-!U�i���dm����d_&����Y\�P����
p�a+M���L�hC�6��D6nD���S>����4 �x ?�;!^���D=�����N
޹	VO������(�n������b��qT�c�L�ʘn�z֍-.
,E�-!ۥ����"^��P'I�1�
 �X�������k���a^c-����.7�C�����nb�W�[o7�!�s>�B�C:��Ga������)�?7�b��?�;�� ��\y:���{eu�ʑ\�9�Tu��g�[E�<h��t꽮�(�N	=�Q��1�[��.C��-��T�t�C�W��5�B��\�3d�������w�Cp�������r'����;�5u�w����u�P�2\�L橊�,|����{||K$�������d�]�1yY}����*��z}��w�%��]��h*�6�a�>��~<��8���]�y�x@�ψr�!�3$-�G�GcۀjJ��J<�}?͘b�!��ӳ�@.9q�%J���g�P��AP��Dl�7D����-�?Kq�k�|����	�-���5��x�;b��٥�!U�ic �Q��.�xT�S�3
�������\����$�Z�5FOR�P���y�w�?�E���ֈ�BU���GV��3�SR®ӄ�b;�s�M�����F��^�5c�@��&'�^��I	 ��'G�z���P�����P?�KP�F��h�V;Q +�:T���+wh�&�r��!��r�R�?sBm<O���|
�P
��h\�=M)�h�Ϭ���P�L��D�&��X ]ސ>��lX��T3hG���m�\0�C>�$�Q]�oJu��O��(�s� ��Q� �����N<FT����sv��o�aJ@�[�~�/�"�h�d������`�dZ�Q]й�f�}���RcxH�{r,��R?KP���	U\4�׫Ӊ��"�eO�.v�u!��0_؆��	��X�MfW�·b�~Lb��V|)��v�a!-p����X�'� |x^^����R�b�����ا��w�tX�qQr�Z�{�aJ�i�\n�*M���E�t���������5��$�5�;�KY.��s����IiХ����,{� -�s���FOa�� �pRŪ��T:�5�J��}"�W��>�����k�����4��/B&P|�����XㅻRvH�07�vM
�De�o,\y���v�8.V���Ґ�ث��(�Xf}=�p.2��g�L��q����*\:��ظ}N�� �aq��Rc��	s-_*��A��D��wW)�˸�7ħ�oޮA*�|ed�(�v�j8gŗ�Nx?��Z��~����q��t���%#��g�vb-ls�H�l��7"�1g�X�S�����cKJ�Ua!����)t���dO@AY�aE�:�[�?<�QH�a-�*�	|J'����������B��te�֙N����lr�
Zh���T,�?���BE��.���ʝ#��	З62�yXt����^1i,����BO���:�렙z����^�'�ߟ'��(��@O�|�4�3^uڛ�)���#�����ݽ���E,
�?N�4���?����]wf�k��D�*�g#�J�X0X{r��E��ts���7m<�ds��ՇG�BlxJ���yeAx���O�N^���P�C���+����1Y;�հF«>z)Kf���s�GM<��IL���?��fg��c�x��qP �o���e�5�0�Qe�� ��j�ҽ��<5~��G75��V�w%�D�HL��)��UN3=/����������*W�0��oCR��_�>�P��>V<`���*hG~�ag>��#�*�W�E�����K�0���Z�ǥ�5�9z��/
��D�:C @:yke��
U��Ǭ���I����!�q����p����6�����` P��Y��Y���|�i7��/������A��u� ,
����z<���贎Z$孃�8��\ ���U�D��i?ӳ1�l�	�Q�m��?���#�w87��)��
0B��75(RP�b����=7��g���n��R�����W��lO�g�?��l�ݒ���n��w��� W�!�O�x�l^z��1�!��FF��5B�����IX�zŴ�Cd���[�}���'�:m8��٬��<�fP8��z�� �Fz0����1jB�#�ap�1#}��stO�~>�.Yb�6���=p۰L�Tmm.i�_�܌Q�@t�6L�YrD~���K2	{��W��o�ZJ�*1�ˀ{/A���\�vp��rv[N��<7���V���g>�
f9����0_\]]]�k{�⨌���j�����0��7H��9�,'�Z��4��(d�f���{:�Z�ds��Y��z�&�u�2�>��А}���0B�\-��D<��ϪY���by�y������Z˶�E�1��lN�Iw��ԥ�y�����ٔ��ԓ>�ɐ=�h��kG�s22�����>Y-��5�ㆳ��듧�+�*����)<�BK���ֆ���`r�����?z�	��?��IiqH�ȅ�X�?k�c��q��v��o��c5A�u7��h�?R�������͵�q�t|����$��W5��.�lG7g>hR�(X�yM'��E���pYo|��
���ro�II���g�1��5�I�~!+%+&I��e�����4���ǣc~�k�`�0�ō�����]'�����nO��K����GZ(܂J��7|ë���:bK.�5�'����p��݉�>�o�)��n��1j�N�eA���R�`�����Ѿ*�+���؟pf�� Q�r�������6��V�����
�����E��_*�A`�#w	��p��.���9¼�*n�����v��0�u�-{���Okz܀h�se�
<C{j7��8ڵ�����QJ�16g~�
��q���a�ss�=�˧d2
	���7���1��X+M�I�Or�s��t]��j���IV#c--]����&�ˠ�SR|k�~̮�O�\Ϙ-;ňЋ,�Isj��1Ȕ���f�M�=U�S:�'���-�@Y�1~���:	��HB�k�r��M(�������Tc4ed:FTe��9Q����d�c���p���$<y�z<b���J����-
����4�dk���*R)���>2,��_G���_�$�5��P��6Z���Q�����ԝ�[���Rt�;�[�~hz��������4��Z͚ߝl��p�V����Qܔ��^8�Li#����ϗ�o� S�e�������2�T���%��pj�o��;��җW7<h�ʍ�K��#l�
�X���4AΝ�LW;m}(�C�/�L7vz�T�= �p���t��
m�)%I���̚����X�B%������/�֌,��˽���OXF�N�#�A�"s ��7���8�g�P��}oq���=��}N�����������[�(=����	�%e�6�1>�x����̽���Mf{i)}^&1�(��-Z��������.o�40���K�-7�+��q��,�rYC����Wk6�u�(��Z�"�儲����p���~�|M�y��Q�:~�ç��n{.��y	�d���
� ݭX�c��vQ�nM�Ԯ��E2 �ݎn��h��*�}7�5ph�Ͽ����2��F��(�s�%��$�[�Y~�����U�(Q�����
Dg�{3�<����7�/�$��Ż���%� 4���\եEE���?�m�~'��(b��'/���ڔnP��l3�\�
��՜�M��\]���'��y�r]52���9��sR_[��G��.5hp�%*�-)}m�P�_�;�3��!*���ԓ�7�v4����n�iy�{n"'�8�����٫Y�4���T����P���rn����Jj6��~�jV�i�B!�� ��{��G���ãRj�����fe��Wف�s����-��ū�,�����{�順<�#��-��|I	��+R���W��"#��:�w+c�xW�<������eш ��B���ݵ)���D�dS't������g#�?�T�z�u{3:)�ݔ%�f8S�vR2���!1��������aη��c�/�k:�X)7gPMe1H܀x�����+�ET��AG�˘z����C`�P{y�� 8�~3.��֑�,ɠq��� �QN:T�M�x��p��H6�hz��^�JJk3L0*^�������l5XO�x���ؑ"~��q�Xi���k�����=u���Ɣ��{�	i���?���;u�߰>��Q�8.	�$EU�ֲ�y�7>�X�Ք�Zjm��Z���N��&���Su���͗�>������r�fc��(�>�0�et�6�du�X#/cR�U�"4���K��jZ;��'�;+�6M�,g^�Aˌ4���Q'ы�Ӈ��җ��Y,�<������=�T�DgK�����+C�����x��Y�q��.�靈�)�q�Y�U)�+�п|}����Ѿ�+���.Vg�ya �J����q��̄sn�r��W���*�rŧ��\��?E��Dal��!a��2>D����D74�/�=_�+w�3�-L�y؇���B�Si�6s��+!{lU�b�$��8���gT?���+�������;p�8�6�v7�r��GR�]y��m�u���4~����%��f�PB�RAؠL��g]I(g����t�l����O���<�l�{HҢa���U�_)��m~:��_c��3�*U d�����Rbu��~ņF/�����ݷ��wܝG; !�l�ޢ��Ϩ���ޝ5�xh���k�2䁊f�nJ�^���'SX$�狍+����8il� ����&�S(���J���.��q�^C�
��U(Ȏg��?��k��n� )AB��9��nT��v>𱬬K滎81X�`��EN���Mt>O�Y�k�#CL�hv�����RH�i�����ٳ�Ww� ����iq�}6�󬝮k��4C��\��$�Iŗ�O����q�"����[1Nc�p6b�N�!�V@#�eu����@8H�ׇ5B�8���9�m Gˈ`��r��(4ߏ�_`Tm{H9�����6�mJ�*��$�řM�Ч(���Ql���Ր���>T&�"�(�@Q�s"��ը�TFW��g��D:۾08�L�e���I���Vr����%!�1��M�������,\A��]�?(ō4�g/�@�� ��͒yǡ���Ln`E�fi�tUw�� �o��<d���_qm�]�>���P�wqɉ�ʲ6~��>�ٷ�I��5�\+�5�7y��#t]��nv�Ihz��A�^q�)�+��[�߆�(��l/]���d�$���{�3���U�ڪm����Ȟ[&��T�D�a��b���M�V�c��:�׿'/�;��l����I�%�~hXAC���Z3,����gz�	r��<$���)J��'Җ��)��]cn<N�@��b�����x�X�N��1`3HPJ5��|M\׿��x�;
7-����l<���ħ�*M���u��{�s�U���3�~���m��ݎP��!�j��d���fH��>s$��q �j����Cs4�>R$~۶0�z���>���d��cK�f�kZ��ٌH7������̸�>�4�$�3������l�S���ܛ�:5�f���������xj���Q"�-��:."@TW���R5XS�XS>��m���4۷�VdK_�����]��/�T0n��|E2e*L�F�V_��b%��=�ks֝��) JmJ�BL�!�y�Y��&���`��E���;�ҡ�9x+hŧᬷ�<s���)}�^a�t�B낺0%��n���M��~B/ٵ�y�]���s�<u97��r�kC��	3�~J%�Vǽ0��;vX�����k<�[ސ:��O�#��F @��'�:���DK���f+�.�������%��u��_���$
�g��S��br�GYRx$z��q��=�1��G�����w㬈5�1�6,Sa�sf�`���<��S�ua��i-�}����^^+�3�.f�|�V�p�	Κ���R�o�e���'1��������	!�8D���Ե��5h4�Bq/��݁���	u��U�:�.C�s!UIͣa�ëK?���a"\ưcFFݡ�Sq����L��a.�&�ж*��B��c:aq�Z#%|Y������=�c��j
�����\�d�(~��as��|K�k��S������{.:^hm}=F��݇�ӧ��OQ�>n�3�i�K��Gى�����ϋ�Oʌ�O�_$�b���8��hh �ȳ.8�GԶP j�=.o��g�yI�=;����W�;�Eg��tnk˦O�͋��B铣��n���+=���bڽ���f�L�ŅW2�gO�o�g]�q�-5��n��T��3.�sx1�u�}17�_�B/�?@f�7��C�o.����A��vԢZ
��޽en�8���/в:�V��kT�:���ݷ�͟Ƴ�;-4�g6���B�M6^͊����94��q6pNfF7���m���BC�І=��AER�A��[��L��t�O�h.��X����c���9��3j�ZGz������:܈�M��Z�ˈ�J�r����ǰ�!��ۭ:�wjj�ՄZ��5�#IR��ClMuɏ3�CA8�}�&�T�o���:$�jц��m�8�>A�1�>]lfs}/b�ȸ�4�`{o$��{�ȈM�Pk�aL_K	�t��u�j��#��w�%�q�!�[��֩蹷��n�}�+������S��Ʊm�G=�%��T�k�W;��WZ�y"��iTg�G>��xo��3��u���o#����#��&K�2*Ç�T>����y���%H|���T����i�>͔���o��C�u��eȧ�qV��訕�/H�C�O��pn��O���|�Q�Dgj<����My����I��C��]�5��Y$.�;O^�PQ�/;������O"Kk�l����#��-�I���uB�)��9@|(_�b�7jy����J�yvs7��Փ�׹96�	�3Yj�����}"����YEWP�K*�)��<�6ġ��.�>�q�g*o4ۥ��/�/����G�:M+/D����Y���+��U���g�P':+�\<${h��U��'%�^�J�Up�|2�w�v�Po	N�߷�*�V�XN��j�g�����+F�g!;���,ʥ[��޾��[m�r�E��$퐼?�Z�r`�&�vOv'����G$�s�Gs�]g��M��у�3UFS��q�''���?�ai�q��̷o���rQ��g�;(��*�T���K�+��� �94#�2�;{����ᮽ�n���CZ�a�J�@=�UI���U�MX��}��b���ؓ"�����׉�''"�oz]D���>�o2��-���nWop�r:�̯!�hX�dB��às�+Eӽ%,�#�#}^�1k�:H��"L����iQc|�fKlv��<��v<��~�`��/��_˥�`o�ד�%iHm���|���v����,��~�(1�\�8�i�I=I��a�7�j���Q
M�;C$os%��b�|K�(W�oY&���'A�+�a��ś5���_��K&����@S����l��Z3��t.A.X��m���#fO� ά�0ؗ6��h:�*~W�P�3a���a#�b�z���Sl%�b/G%�!��%6��\�9'������Y��ڐO[b�l笌�P4dMY����Q�^�H��5)��T)7��"��pT�K7-�z������c����r��择�R��5�ڨ֐�)�W"-���v�˧i�e�E
T?�	O�Ο��@ݯ����J�[�M�?�:�:�(V�y��Бj��F�2�5
�J&JW�X$�#��e�����j��0��R���bΟ��]%�P�@�]G%쩒ߥ#m�J�]
"�\�?n<�����b����#o�0��L�8�I�ӣ��9e��|�F�+�!1h�p@�K���MD���G��/K����˛�^���4M30�H�xQ(��ˢv�"[��� ����dt����L�LM닞�f���Q(m��5�=�I%�H���B�~���ɮc�$�C����Va���V�J��k���m<ļ��|q�N�%L/���S�"L�q&�
��0R�O�Vff��P7�����LY'Qc��#����oDmO� -W�zi6FM�X�hp�uĉ�G4*Ku��Fc�5�Ø�`c�"��2ܮT7��Ш�Z�|^�x�3�,��a�п���>l/��T7IM�Z��K��6z��8F����[E*"d�`���a ѽ�*;�2��dz�dQܲτ\n<%'͂ͮ6�3����}�jq;��=	�UC*N���^�3�4��T�ҥ��{�f���M�9�9����N������'���m��Ό�����!�3�_�����^�d&��@��Q��S��M�,A��'n(�V��=�O�DY��R���5�խj=�K8s��+��;(�8)qۍ��C��s�F`�p�w�*X�s��5��'eg�RX�{h�0c��BQ�`�A	ApA����eQKk�^�*E���~�:N��=Ĳ[���a�է"{h��{}�~�?��J6�����L��h��Y�4e��8�oQ0)J�y ��<aX�/��+/b��#�ѵ�o��\j�L����K`b�#T"Y�^�G���� ��b�nD����ee�YD4S�3/¾Ȧ�j�.RH�kx�e�e���!�W�}!c&%���6�Y�Co��u�d�!��Z�H����MF�j����@��M�GY�Յ7@����Rc�R�(1�����)a�·"i�u�����h4]_��I���}�Rx~M���"Ɵ�����_}Q|u�Y �� ^�o�?�T<�F���E�����i*1�`B!Ɯ�4�b��N�j���!*�	�d��A'��q��LD�x�ŀ�b�	xL��֓��;� 1�%Yb�C0Mwo� 63�{]Y�n�wx��"�ej�xԙ�j�X��9��߱>����Hp�ol���*(ߎ�1�U 	'��YCc5��à��﫿�[�S-���J�5�MLO��L�K�q0��Po[�R"���M�����f`~�Cu[%,�6@��|����J8��ę�\Z���f��<n=�u�q����}5[�,~&z��{����;��[���늷����>�\r6O0�=�ػ~��%菍]T#��E�}�@���
ć�iZ����3V��m��';�,>\�u3�5�ر�zU����IS>�\���%x9�uezk���������u�D��G����w|�Pp+�	CJ��5�,!�Pe��P��T`e/��(�j�7��=�L_k�F;��XҌ�$/������τ�b�[017��M1掩$�m����khT9����t���%�a����W�t�g�u�k.WW$��ِDDD�&O��hpq�=�Hb�*ڞ��Q��] Eo;<��Pd��Ej	o���p���z[��_�*.�:!y�X�P܅7/�:V����B�0Sv���,N�&,����/�n��(�V�����/F���[���覡#��K1���I����4�����Al �i��ڻ�Ƹ��`_j�Oe�A�@f��xV�-E Td�nbsH;`�O���W��U� ��iG�����>%�����������o$�7.�?�(�fZ
���A��|��|�l='D��'��si����r�b
A�*��}��Ĳ�i��2����_ְG+�ҩ�qrJ1}�D�v��P��A��lz�FI~�?�M��?���g��7�!O:?�#�q��L�&+������/�	��/�rA��c�u@%�I�y �z���� �؄�חMW�ui�w2�1�!��}�%�$�	V)aZYT�@�L�	wR"�
3����}��8�]���������C�^�\y�k����@��{���j�a\�3��ҕ�;���TP{q��`����`_�S�'���2�[&,B��{�`�ǈA�x?�j{^	�j��</t\Qg�.�k������!Y�����
�y���d�inn����a�Ts�����~Di�X����u4�Ù��&���>�	ɆN���;Q<-&պ��3S`�\8�d�`"Q��-]�B,7��7(E�p�dZ?�%���#����Է��Cu���~�*׃/y���|ow��_@��lz�N�U��H�/�k��ޑ%�5<ΒM�PG���~n�T$l��������)�Q�B����`��];i���Y)�S�yh.Um�pc~EB���̭����=D��Ue�2u8V����>��>Wg�B��Ǐ�|'����aƙ�z�V5;�e��!�)�1R=$�-�:AH?\��4Lr�5���u9��o��Q���I��߫\��LKF=t"�Y��a���z�sZ0�l�?v���]�͗�<<1K4�SV3���������@��`NX�@��K�ju=��Q���h�����x��4��Ii3�W�s��b+��vҠ	\�{b+H^�%.nF�&Q�|��H��h�O.�!�
�n����,��ʍP��k>��#�����T8���_�կ�'{/yx�z!@O	%��K��:(�Y;�_P���ء���Uw��i�R*G~�M����v^�d��f"x(~c�ٖ�a�l�Ϯ�1�pjM�ן��A<�)p	�`|�;����!OB2��r����Sp��޷?͈�ׅ��YE��{)2�	AҤ<[�5�4���D^=�e>�E�`)z�mEg���Z
�vxU�� {-4��f�|��x��o�/TH�	�}�_���ݠ&����}���y�h���������I�,��a���"�/E�i>Z�����6?6�ƪ3������`�� �#�X�$jW���,��D8��c@p�]�%3XU�G{� K�_�� e6��JIO8�Y�o^j��Rjf���͟R�]�p�;���w�>֌�)�a�u��x�u��n �qg�tJ��/������������>D+�-��h1nyʴ�]�����q��Yi66h��ډ�w&��]�<A�*3�^O� �V�������%L"�ٌ̤�i�� 7�+Z&M�#�j�7.���js�g��0��2�|bs����z���,e4Y�!���AHP��m@{.+�xE&�h$Hl��>�H��u9"�[���nDS�쏥^��a�P~Z\u#���*FIZΫBH*���Y���W�!3��2��aJ��F�I0_}OY6��Lb�H�s7��-�j\�c�(m�n#�Ϋ�O4K"&F;��@mT����������]�.[=�
z��w��p�-o���ۛ[=t�Fv�"��4���p�v����0�Gʈ������d�a��|��r�5��:f�?�ḵ�7�3����3B<���v70�Ԓ��S)�笂����g+o�ZSs��p��ˀunF3=i��U���Ѿ�O� �f}�r'�f$�"���N�\p�yk;�ܾ7�œa�b)&�v�(�E,�W)��iF>��\�'GUQ����#�J������w�粜(`����Y��ţ�$VǳP�3}Ed��R�c�]�}_���b�`.���;Â)AW0��_��q�����)Q�0^_w���,J1�i�/��%~-�oqPK1ց�:w�o����A��e)��<�C��vs��`I\T6���>��Q}�B�`w�F�'�N��������m>�%y-EJ�1|��v�͞�n��������r����]�����^��0iN�b�X��g�4A6R,�JLN�N���S=$�3��aKh�.T8����xTz�9�LIQWhU��0��&�l�六�(������4q��ɶ'+��6͍�����ht�6�)��W��|���4���&�5N�:���{}VhE�j#$��W�@����Fԩ��E1m�r9�poc�����Ƌ�E��8�L�&�AUl�����?�?��Hc/XOƸ�S������"����0X�Kmd�L��]���V��"��{�̻��:Ȱ8��?Uzn�!B��)���h&�H8*���ì��:}�%�0T} %WS��q!	?Y��+kIe�0���-[3�v���m�S;�+�\����㿐 v�3P�9���Ƅ���Q5"��a(4���@�00�\+�~��aN����4�Ck�i�������.��w����[���D�=��Tǝ��=6�8����3��$��PC���L%9|�Q/��U���Q)��m�E*)f�;H��9��Ѻ���q��Ј*W���m���Ҽx̲� X��OJ��*��4�sr�D����"��G2��-���(�\��j�d.'���n����24g��$wz��9]f=��
��D��܅	$܁%�8s��	�,�v�V����5��0%�c��T+��ˑ�*ʏ:a�ēz:@v�n^���e���i��)xD5�Ҟ�c�)�U��+��j�<�˛�Y��N]4��Zp�Ӆ�&�F��<Ț
� �!ob'HCX���UM��y�H��}�O��-���}]� ��3A���(�7���p3�g=\B��<_f�r¨��ߟ�b#[В��+`Ϝ���E��F�������i�}�٬�A[L�}���RU�E������UU%�|�E=�?������t�4� '��@��0�N.��P,�Hz�b�g�y��Ӈ⡃�D,���3�ѳ��t[���y�-nQ̪�&�������qe$X�F�Ϻ#��ka��r�)I�c��� G$��t����$�����eӗ����
f�B���*At�l��A22�Y,y=��d�Ǵ�:7�7��8���Fg/�q����|q�5�C��	���EE`��ק@q]�V��"�b��]�&��m,D� ����\�8[\T�u�M�Dx�����x�OF�쑣s��b?���Q��H��O�F���_�Mp��ȁ���b�
�^ws�]���y��K`F�ˋ���bG�'CI���	�1CA�`=D:��p)���Vɇi!XY�#7+'�R��a"�w��3E�	p� WA0���YM����k�xfl;?\�@�bY1�=!�#e��|��Ҹ`%�5���UU�������Vw��f�D�P�T4��gl'Lڣ$ @��ԟ%��O��z_=!��R=X�hfuE�{���L(C(�/���-�NY0��넱�GL?�� V�� @��T3?H���""&�3�}Rz�.$��P����8���a�?G5�$��=�*��)ci���K��nE��s�Lc���M�ipjg�v�b�~�`%��/�~�t�&v1��5%�/QG�,4�$$�s�ݲc`-�Тy� "f���o�%\��y ��N�A ���c^2��l%�@�}��\� �D4��K�Cx�)|&�oVH:Ha�M�9�]ya�F�	y�]v0�=��v�`&�W#ε�Y�o�_Y�3I���\Egk�.�tg&JЖ\b�&A���L�/�̔?X��B.b�*�>�+��)�3=����@��������n�a���'��ǿ�kՂ��d��é\��Z�Ѽ_�DH�^`�
c�;Ą/�����rP�}D��J5���&���F���f>��j�6���g�3���HI����X%}�D'Y � �w�O=O1EY�f]�����Z����	�>%�m..�xU9c!r;�~���}�ֻ�C��~\�x�z���P�� 	�(�x1�B��Qe�ok���4�u��0��x��	��}�:LZ��Ѫe� �$��]ׁ�_DU�F�M?S����v]E�?�"�OQM�_�	`m���a�AV�,
L��`9&�0�͓C�=�}��x;�M7�Y�9��)�Gaz����çcK�?�+&�L^�H�Evʃ2a�cLxy)�Ƭp�����~�w^h�+"ꓫ�i ڟ��w�%�;�[�����N{n��<	�/ޙ�e��y3���|Ö��Vq��a-d ��8��j9�R2q���"x��Ӫ_�?W�<�0Cx�2J���]:*�#=Z�S���@�9���~��r�w��Ѱ�MpwwG������W�z�Jo�BC��5���ш�oo��c���' X	�_LU��t�B�n)���k/���#�z�$So�XYW�}n�	�u�^"zʻ���}~A��:����,���;�C��j�e@H^����T� ���[��y���k?����v�~ņߘ�F����Z�z"~�618�!jF�.��~M��eƍ(���~#�ᤲ��[l��x���t�%�ϵ=o��X�r� ��K3� �-Ӱ7U�,��+�j�|�`��ͶI3�8�k�V�EǇwv0��ٷb��6q0�~���g�՝�������dif� <ؠ1v�2�[���}΍�Ŗ��o;2��p�"a�!�~v���t�3�"�f����ۛ��IXyPm���2܏������ ?;B�y�G�l�X,pR���4�����Pg�~�3� }�]�DsOx�'��O[[
EO�79�hگ�h���m? B�R�l�z���	@%�(U��%�&��/zE�Уv�7���x��>U������ޑ7�2oѮe��-��B�s��D�)�[�P�����w��!XQM��N�ͬ��2qje:+�gZ��8���2� g�p��"�P4t�_�}YJ� �
�b٩*��}�6 ����<Y��K������Ȏ���]b|7�r7�"��kk�e�g�a\�#��ҁuȗ%6��� �z�2�/�y~��o����&B�4t�������4
��`%�m/�GB�o+�|9HLlN�LV�P����>R�&J���V�?�@�`M��'�c���TK�V�����xi�X�섳��c����cF�p��A�e�-ю�TND7X� �?�+C�?��"Z�#j��W�Pq�n&���� DhH�ْ�0͞r����!U̮��Q��Į
��+'�;/B .@��&+�22�3��iB�������iN���Vd�3Ɉ�|�@Xn�YC%�h�9
���]"�Ñ �J����r-��0�r#Tq��Zp �&��Ed��s���i�ۉ�W�R��|FW� �9Y�ybJ��3L$��d��0
E����t�1e~�c�jw���!-(�ݒ��p7����-����-{��a�?O}��gyeh>[(�*,�ۏۖl�5
�� R+����e^�c�<�7��?��ȋ kQwʬ#�ܳ�g��hYݥ/�uS{�rP� �G�(R��L㧁�X�q�n�	9K�?�aV�ç��#ݘ���Hi���~�P�� D5�C_�c���E}V�Yd���y���{��}��n�H�7C3�-��UF}΢�9C1-	r�j������C�A�^��`�
E�R������ߤ`���X���%M@��%��� �k�>�_����
~���e	���p�]>���t��cՂQ���T�J����h�C��q?(�X�[�%�t�4n����M@E���C��r�_�-��	����h<�]�Ӛ\)���m�Y��B����j�a;B(Q�Hb�{��ŽZR��A����>��7�7]���a�/`[g�i�_���*Z��@������}�XX�z�s~�'��S�S6yaa�$��ODzV������ɒ��D���啰�B�zR�i���	t���h����A������F�� Z�K�a9�B��h�`�1=J=eN��ޒ�H����в���ٵ��3�Г۱�ݥ}S�PQ��i�	��1��H�*�ި׾���r^�ֹ�P����!Y�Z2����Y���c��h���!��}:�$"Q��o�o�r��=�HUH���N s�Mӗ'�8�^�)s���_��>�Ve�@�2|B���
6��UH��@&�*,��t���w�4qn��JK2#�����FQ89tԵ*"���`[]�+�N�3�`\|��}��>�8ի�8�U�"�I'i�>@�����_1F�1Zlr8P�a��9��K�d��jX��YZ]P<b;o�^��x���,**�,Q���f���f�R��{���a��F*%e�itT'���{��m/U��H72���;RɤV���C{���<90��n�S6�����L���ZTWVP^��˅?�ЌU�?rJ�e�Fl��h�;:�4AꩤaM�52f�g�'F�ܺ�yZ����Sksf�K�vޫ�6��0;��OF�md3@�_�M�Z�o�9����?�[�\��b[ے���uq23N ��+�@Ge2�U�jo6�zp���вxH U�IX�O������������CI5��͋~zm$�y�s�g�)C-�D-��9���Zv�!7P�`���07,&L{���^�J��0gֻO�������d!�&�N��$��?���]�$�;'��)��VX��*�=@y1(w0������l�NS�^�n$k�-F���	�.&����T�M���}���i��;�{<E��ҥ����t���f�D��J�^�A�,�[D7;�
e{�P��[n����Ր�c�xnNpKC+�H�6f��~��~J��i4�[��*����6�]G�(��'vI��|��kq��2
q�����I����.q辬	��a�[T������������NN";1�_����q?��+�(9��м�@�HK5��=�b?�5���t�ᡱ�b������}���e��'f�Rݼ��A} �� �Q��Y,��ь��W�N*�
Gp֌4ߑ9~�&v��2*���{ ��������	��wgpw��n���n�!����w�:���Uջ���kvV���I�����)����rr������ͅ�V����^bcT�폃����d�/��y.�,V��Ү�v��.�s�+�Ot�&�b"�4w{�-�X9��u����M���i��1�-���j��Q�QP�F�HJ���%A�C[�veՃ-tY���V�#RT.oK��d�ƺ���N�?��d�q�S���
��3rtBl]Nn	h<갯��L�������/���-���I�wW,������~7O�d���h�5�҄x�����Pcn�k]���w����l�"���}}�s)w��]���p�P`b�L�s7-^� {3��g~�{Yƃw�LP����i$�+x���$���gsG�ד� bh|m,�>��ʔ:��L�M��*YEj�Sˣ�����ȸCo�4J4(f�?���4��2������K���V���O�?�xy���ù�Bȼ�ĵ���C-4��#�Ȟ��&9(/�$�����]�_�6A���؛'Y�0?�s�����e�Ҹi�ۻO��y����VK�m��zX����������ow`��g��V���i_�y����7�!� �w�vT-��fl�+`g��Յ�����Bt׌�̲�B-!+�,	�!*�^���0�&J/[N�#F�&����y�]g�<	"|������Ŋۧ�&D1daxI���¿('s)ڛ�D�,�����H���"����D���@o��R%���cJ�#G�n0K;�f� y2�A�u#_a��o�� O�6�!�+/کKQ��}#VX~N���i �������D@��h�x�ӕ�p3�W�mf^�.�����jc�ӯ�	݉7!��*[ɾ�*v��`�fA�q�jY*��W�aJ�y�Y߉U1X�rG����K>��JZ��3i�d%/%�M�YTi��ԑ��K0�+.����m�PcA����8��ٴI��k�Ԁ��lQ@��'|dY�%C��L�v�b
��p	�+B}S��>pP����Ѵ�������G2mL��PK�Z\p�Y�RC�,���r`�D3�����v9��y;Hͫ��<`"�PQ?g,B+TW꺼�����@�d��;*w8���P�0�I	'y��6�O�ӯ���8���L�"a�o_$F.|{fB��W�<vn��_���Z�Q����;
q٠�ޅ��1�c��7�:�kF@�T�w�'-C��0cJA����DH(��D�}1���t�B�vN��n�(=� �=Ε���5��L�EMIȒ�O(��5K1d��*���1����Y�C����JcmQ<�6��Y����=��c�1=��-(
���>R<5�/́K���vq��(wbؙK�đ����` ���/cfU�W������6JA\k|�� �G�kXlLcW�e�A���킽�Im3��5���a�7B����O0Q�1�Tf���If���ڒ�P^~o]8��G]Z ��i��/�����鄃�c�w`+4����'5�B�h�h�7�.f�[�����	���/�cO֠c�������g$&!$(�㪛�(?��2�u�B�,bI�:��=M�\�h�;վ����[-9T�;�Q������T]�����خ�����d��k=�c�!\J<�(���X��V�@�E�����VF��0p�X)��C[��Ì߈s����R��T�Ԃ���E0!�`�w�8紉p���?�4��E��s<a]�1��%t8�0�hz��q��� m4�Ꮽp��;�׫��Z��E��̖~Ibn��0k�T�p/7��y��O��.1;=\C5����;�$�,�|�w���w솃�<���Fɉ��
W=�ܥ�@K��(�8=p������Ø�4�ȭA��@H��&"/m���3v!	�~ϔ��5"�_v�?�98�wh�Ί)5�f�9�/R�4q_�g�IE�g#?@����B���r&���^퀅�V܋��P��'����#y_�Ξ^����;��_6	�^�B��P��̂�@�Շ���y� Tn3i�2Fy�.� �~�ʑ�+�Cmf.�����ڙ�A���z{)n7S$̸�E:�vp\≮-H���r^Mc���@*���g�NHN�U1�4�-vr��<�i�Eu��� �ݱ�H'��\�	;_FD|�d%�����PC߉�\еq)�L�N�?(ʮނ"b���J��D{K����S���'�tψW������<����Lb�n���G��¨@]C��\zrH��Dʭ��#�˒�4-/��D&3X�1����3�d� �������(!-?����������߲�B.���0�3_ 	�S�΋ ͧ�b�4t��HՃ��$�$�>�SyI
��^) %(O|0��֨��DL?8(;ͼD��~iA�,~��D��ג(��t��qc�N�BOc�������!�7K����q���z�y"���ӫ���Th���cJ,���&���91v.���Y\�2g�R}�\G����:�����S�NC�;���x��;0]�H4��=�26N���*��ӭ�,�((�"�c�f}|.-������T�H�8�����_�$�E����I�g��(��`���9�Hk�QE�\�~םf�;�� ��0Q3\zړ��O�Xd~�cȢ���[o�74z��t�O:�,�?��������k��$TH_g+J�l4�#��[�������B8�+
��z��bB�p�3���%-n]��*B��v�� �3~��:�M�!�����v/��ؘ	B`fD�c�������<4��aܤ��¤""c�- ��шOU��~�1�Ǒ_A����"�4;�t�9��ֺ��s�'G v,o'�K�z@ ��̌�F�=b���jZP�1�0I�0b����[Io�U�|�Q�;�R"8�E݄=ͫ.�������zl��>�_i|(	�@��5���	"wJ�m�]g��	��_�EЦ�D�M��5K�f�P<�E��D!l,�jE�@7�� �=C��i�?��eJD$�K��j�l������V��SD���Ɇ�А�� ��_C�8Y�w���z�H���k��k��+A����J V@
 8$WT�iB��
6_1?:�z?C�����(�tnT&~P�~Fܔ��J?l\�*�X\�_%n�f�x��b��L���.(��[8W�^
�ߟDɧp�*���g黔/�5���};bT9[��荄頻F�2T��#"@���i��"��8ʄ��#@��H�xw�,��	j��
�,8S((�����Ǯ��(��Y-��[�-4˕�`��5*[Q֨\��ۤ�3�+jsPs���I)�2䠿�DFRP�\<K���@�	0H��L�{G��Q}�Nӆ�Gw��{�0p~�a�ɢe���m�&��&ȠH"u*�mޞa4C���!Ľ�\�����ͻ��g�g�B���3��xdc�0I�<�TΝ��v���MwyW,,�f3V�^�a1���#�l�~�a�B�trϪ�`aq�a�����	p��b�TR� =쎽���R�=S�F?>8fSCe��w�(���o
��;}�!X�C|�
�@��^:J����	�w@R�$��[�E�Wp}�lظٵ�3�#t�#���@����0��԰��r*���ExB��Z%�&�����][�a�8�:�J��'���ç��G�M9����7T��r��[L����B��	I`��!u�
���SI���s\J�2��A�5�<�e���
���b�T{�LU�����k�2���#B���NZ�4�ڵ������!�N:ʋP ��uoVd���q���yb�G�>��@��T�A�t�J�^�O%�"O0|hȀ�6���7D������������h�IS�}>P�,���捻�Z&�@�6��=��R��c�q�4�Q9R�<{v��!��ֽ�U�����X��bx5LZA1l
���S@%Y���j9̚�r5L2y3�T�n�=\���c��/��_~Rt��	��i���uN}�/�rh1#uNBs�=��SL�Sӝ�?���~.^m�g�8��n���KP�*/�9�TG��|�H�����G���.��g�V����[���5Yk��G���]�u�V�uC�����V�CF	>:�. u�����B���~#P3�o���F�q���o�в��&���q�5���� �-����E���ӂ\����X]Su������i_��� �9��_��E)o?n������<9�����"�`h̏	�.����b<�9�c<�{�	��2*�_O��Y� ���#��K�	�5��%I*իl��U\[r$�����|�<n��42\�2�1�փ�]{O�j[_N�]í�"	:'R��!Zll�U���%�����䯟�F&�fJ�[ٔUX�yڪ��^1d�1j<D.h�B�b�Z������Y�D��f�x����i��;��E4.����}�q�u���G��<�l�P�"��fOzL���թ�9-�w���=��"'k.cM}���W������-+Ŵ�����4�" �!?��:��jd��s��Lj�0��E�E�2�m��u�C~�j4����Q��J��Wj��[ޥ)�e�Ϩ�WAu3�
.-{oZ%��mjOU�5�ېv��M6^J�tQ"���h�K���L�ދ��<2n��OoC��n����\�0 ב&�@ll7T�xl��@l�/�i��T���6L� ����c0����е~��a�s�y{U?�5�sQ�V
J0��[mzz�'�	q쀈F�+d^��O�v�ǶhI��.2����).��Q���ɕ��4�?��*���JC^���_U@��}�_�'�ӸSe�����yk�{�6b�O/��y��
�%;�E/�vW�e~[7��Vss*W���#{���qMe�J3}!Bq��ڶ]	�p���z����Q~��d��1qM�Utq��w�rKm߾��XT�Z�iD�e����~�L>`�'��*i�UUS�J��o'�xB����o3-�h���ul���u���~�:�x�W�$��vH�D*ge��^es�nթ��9(/�je=S�YN������;�+��.h\x�%������C�Kd�	Y?;�^�l(q�D.��z��5�}.T�1��M��{���gd	b�I7�{���|�yO��kԲE���y���������sB	,f�ؕ�� ��_���M��5k�+]/sT�Ly�7d�N�{�,1&g�x?�:��:�f�F?c��z�G!�-p�w�`�~�V������Y��#�]���!FT�#O0�^c~J$U��_Z�7r]=%��ź�:	D�+¼����lj�.��]�,�H����88i�N~��n	
ڔꀘ�BL��7z}��w����@g��5#ܼ�wg�s/��H��c3���^)��4t�wj�8���V߁S}�ְ)@g�oZg!A���hCk{wB�%����\��E�y��<]s�����"k#3���m�"ͬR|/�-EZ1�H��>籟��q|���i�7�RZ%H�~����q�����ۜ���'�?@R�3nW��o�d�-����6n�las�g����ٔ���:��ϭ��UoN[9z?��Nbu5�۫in�?��Z���Ģ|/�+��W�-?�A�yI �� �{��k���Q��fc�/��^w����4�Ճ�j",��Jęb��gg�%��o�Y7d�Ųխ��1GG
L�[����abK�U)*�m�s�GI�k;���N[,��e�j-?��G�w��h�?Վ|��T7;�;bd];�8Py�c[�qL�ƶ���"���xB�N��q���NR,k��m�>��wR%wN��<�1��ZS���N�,q@M�wva!d�Δv�Y���-e��\s!�Ẓ�	!��Zj��5`ݽ:NNX��Ij�̖��*�x��ᠷr��qd����]
��ATiy�~^���{�*��ǒ>�����b~�)8��[�	U�+��Mr&�^:aI�.m`�X/�_g��z�QX��;x�+N֭+����D�׫p_`-�
W-[�q��z�E%�g53ط�x>x�G���^��{��h�ǟ�����q
���F�8����'~��PՕ}H���Y@����K���9�mJ|�����s�	?ιL�{�j�r����)`��CY�<7BYk^ͺJ��K�C�Y��p��
�����k��VS^8!��������7�,A�g�1��T���J�f��0X�I�)L8�m�Ӱb���t'	#%2TlK�^����&�V��޶+�~�|��rOA�y	,:��r��p�?���=�H=�	�}Uo<��}��S<i|ئ7���u=7Ki]B��U�7I��+��q��4��e�Ϗ����u�-SE���0��K��=�K��u8���һ��.���z7Pǻ�Z~�&��φ�������:�H��dq�M����G�-k��Cwk��A��� ���?�k�hD��:��j�����n�I�=��{���>��Ѭ������ᎧG��^kڱR�nM�	o���dP1W���:��r�1��N��������_�w�����ޞ�i^W��~�\
�c��8�귦�"_D��y�P$��S��^:)ߒV���I>��|��[����$	=Ԯ���Kk� ~]9v�	K[A��M"��`?����b���_�|Z��7��	I��С�[�{�6��_����w�j�����^>��躞(���H��{ `�س7
����{P��t)�o_/��/e��=y�g�ή>W���M|�y��G0����I`�J�Du��G��0]�7���!�,���F����uq�;�����V�:j��;2�u\/��� 3�f:B!:���F7P_^��Up m5Ӂ��V뵥�e�H����������i�	���H>��1bx�Qb������d)�\�.&ޖ�h����H	�op٣J�u�;�z�_��z�b���W9��
��?���q�bEO��O��]��W`����fC��Ċ��G����n�<��zF��4�Ua$Q0Ӱ�E�d?�ǲ�'�g�wc&vV�$��P�Gƴ�o��V�ٟ`����FS��".�	F1����m�~�(�"�(V���h�9P���g{G��Q���n@�m�&�+rt\]ƃ�j�0��kC�>Imٿ�ux`�E��_��-�Uo���`�yL��^��5���JV��5�,�����v������N.�n�3@����N���u�+��>k'��͐�t�� �����S]x݆ϡL��e����3���S�u��2��c�V��G��2B�������b���1��$����	ß
G�u:͍>S�g�a|��0;���j;i5�E�q��^� E;�W�&+:�6s�)BCc|����VR�h��W�������C�O�ц\����EW�ª6��i�k͖c���py!z��rj�$GhF�O%%���A2a��[�Ā�ծ�3pH�iM�����۵����3�@�8���\�����Sypu�.:�\pk���F��LαF�Eh�AP��x���ɗ:u&䡬�zu��ۆu�ԫ;��q��u�������2*)i@���2Zq�nAZ"������1@*K6��g����S��ֵԵ�̆�b���t� I��{�у�$�O�ޮ�[o��׹ɰ��^��a"�@)�~�Yb)=�Sa��[�@eO�&v�f��Z·�?�c��&���c]��d~��<����N�#C�/�- �C�y�.I�aV���J'�U�������0{�l���|<G����*���O�de,Mڀl��-�Szj�~꾻��"���]��f�>7h�^��@sV���� �%��cA�Bյr�g��a��d�7x�O���'�~x����o�h�шUE�;`D��e���$���)�ޕ�{�GY}et�U�-Ͱ�;v���@�0z�ǃ�<���Fndsq+�#{�/�Ӣ~�SuI;&�Nj9U�_;��)�1<�i287�u��c�4�H)Rv@@x؊M6'�2���kj?��e/T��1�U�Ts&�8K@os�ٚm�����E��bxK��Y�|>gK�8�-���!m
�]�bI����-��D�k�a����S=)kH��u��]ĥ�3L �|2���(h�wm�@�r�7�qUu�@�?ߜ�#���+:g�ʻޔa��g���ѧ� �H��!O�JO�.��$N���R6���4�ނ%L촘p�G�d����nf��׊��K����K:���6��KVҶ����#�9��m� hC�ǧ}O���޶�����V�M���&�m�o��|���]3��_�V�L.�h���<9XPz���Qk_�(I�E���d)#�7JB��a�V;���o5iJ���^�5��&��	�O��
;�2�1��s\�<R
ۛ���n�t��S�^&`V�'�P����}��P���7���i��sR*��*r[/#s��¨�%a���X��i�f�Ld�4��B~�bĬ\�p��1C�^|��.�iA,5�U�Xz��{8�쉋R�!tN���3�I��a����v|w����q7��]�ЍH���ZԮ�*��N_O���%w7���h8�]����H�tm��!nCe�˹p�u%��I�Hr��`����r�3 ���I����D,.�/G���l�]un ��6��"/[��
 �{p��Y�LF�_+b��h���Ӂ`����%��ѕ�)���;��x�o���_u����G]�~A��as>�=�2�4�?i�;[��p����O���|�Osu�<N ��Q��lsKHJ�h�����|}�:�z,��Cms��[p%v	m*!�;��J2y�m��ϧ}�	H�������rL��|�{ ��\�7Il3~�Vr?cL�U]��a�3<g����ޝv����yq�
�̨
�e=X+V`��o3s�� �ڤ<o��;Y�i;U8U���,�����>��	��~�����F|��Q�wl����v�����JM`����#g���MT�舶���$j��1΅���I
Git���m����~̚:�#ce�)�c�8�[)�!�9�s"Z�r�?o��68T���s�,?���3�R�����i�e��Liao/S��@.�KB�?���Fߏ�L���$ɓ�WІ�6"#��m<���XZ�:<�cy+���P�x�(��	���G���������3��}:XX�7i���b�f70�+����)��W�FZ��t��1���f���[mEF�@��zr~����:���h���?��KJ�C	bu�6w&JrGJ+�~։�_-���(@��nR�
��k_��s��e~6ĭ�A��e��*�6V���bS�	a|�Cە����0�ߗ�oz���[�����p��e��zw�/��6��W�����9�a�&OC�S���1%a�3Y���}<�M�׮��'a.��&�M���T|��-v��Y�3�]8�.9T�5���Jjly5��h����]��UטƓI�jL�{N@�Fԋ<��s��Ф|x�6����VQ_2%+��[��yBס�3a	�u���4KSo�R-w!CQ��%��c���ޕ�����*P�����"Z`F�V�]����΋�8�g���Eﻔs��Z��m���kd���~z�9E��㰂�Aь�H�����6�12�q������L�Zl�W���z�q��9�����J�?�/��r��z���?()�ЎA��1����k����	���i�Z��1�@� ,�k&&$�cl丫��/�V�-�k�;^��6���ϰ�V�U򶺒N7	WMGE����׳�ӦN�NHIe�HXe,B�/.��
�?  S�@��z{X3��p�[VDg�@��������R������Nt�p|��a�~�����!���^���ު{�X2-�G{^�Kh}ܞ%g�W�V]�yM����(l�D(�W�[_م��;�\���+	V��@�D�M��.˲���$�ie���,��d�ĚH�P4]�wwz�̐}�7���.|;�,�/�s�"	
����&ps�5R���,>�,h�wU�E��4��I!���)V�~|�J_��c�N
gYz�2軯�J^��(�R�lGf���i�ٜ��c`�l�9̚�"�
|<��?p#d�~������f��3 `B�k	P�gI�����<��n�������m�9�Pۗ��L��}�
}�bZc�~�s&���j7�b�O���e�D�9hmh�K���*����&n`8��2���x�������2�И��з6<3=7(d��i��2슜���z��g�ղ�ԎʾC���/q��}��a�c^q۬\���p߻� ��=Mz���i	=�#��p�LhƫP��u1kF/��y��t�Ml:��gcEI��E>�#���
��6�(���S1!��V�j����M���6V�Nذ�Ede��4_��&\�X�����4��������򢋏��E�n'���k��;�����e�Z��
P7qlAQg���w�ek�!c$'�Zj	(٤�6:���W]��"�G
8,�3C��Mz(y9*��$��C��&*�i��_����a�T7��'o�:z���ײ�'�Jk[�\��~�h�q�j�Pd�i�5���=́�&�2q�<�����_?�� ��*xx���KH�i�a��!��X��ϡn1�����c�6�@���hw����;�m�|�_=?g���*:��c9�L����4i���2����ۜ=�2�ݫ��n	Y�=|��pm�A�,�($-���Ƥ���l��X�X�E��%Ȣ(iV�i@���6,R��6U^�Lx�y^\vmU__�q�JP�\�ѿ����>)Ѹ��Yud���Xn�ota,�b٫p���ԑ�@c���4�I��p��يA�T��ǵ1|m�8�8w_��И	��A�q��=d%�q��ZU��u�T�+.1<�r��=���be6:i��T�p���M�Ⓑ��kȁ[qq���y(:�統9e^�v��a^�'���k�~J��n��ɮbM�C`�a`>cTRmB\O��B�V��������R�����T�c:�ƫ�Z�eT�00v_i{T��5p&��n�C���'���K�6��)ZX\��v�.S|$�C	�p}�P�9(�3W�[%�� ��Z��U��!emm]�SK��"�p06϶C�\�V�Ev������E�֡��|���~����ԣO������)��
� ��hU>2���ړR�"��e:Ā��r-y�S���-�M�*��bA�^����������E�O�N"żo���|jG�df���agr�+��T��,��ء'xP� �����Y�p�Vc�K���uW_|7f��BF���d:��G�N!�Mk��\G�����1�{��dG��dW9�W{�����)��3�Zʖ���ŋ�E��/ߞ�뙳�,x1pG,�������y�8¨���_@�.� �}�(1��V0C㝹~�?����v�����l�?Q������g��5A���Xzb�4�^�����Zu��"��6�� f�t�)��G����'dכ�j������ؤ.��;ے!�4�0i�d �s$�~��&l?v�D61zŸ¢����$cck�+���tRz0��Y�}����& jZ����@Q3,����u�������������;�O�:���&�0g�-p��3 �(/b_�n�z�_۶�SLTX�����_�;���&�>��酃��u�iX���xwC�<[a�Ev��ʀ{���9I>(֍���{�,��?V�}�z��6A���v���$�G����V	�%A�'(�� ��=�=�|�?���u��#�dW��Z���.�1��d���AԤ>�.:1�C�R^?�����+�?��U�����h+DE�G.��[F���>FG������~�b-�-
�O[� �slV�&����+����&& �� =��&%d�v�U<�=W�� ����D���PC��mT#(8��3P��e�B�>�6cDh��
���$�Q��/`�(��}�"Tn�:)��8'OZ�˴-"2ݷ��${M-"�����Ya���WB� �� @5�z[e��c�
A���U���i��r�;t������.۷0��ʑ��Ѱ�����]�+)+-_|x`-����u
������UM��D֒�������5|��G�-�>��[ќ�i�Pd^�|�JFfs���-4��V�C�:�@�f�Gy�^[D=�c�w�>��v3>f#z#��T�v>�ɩ$t�Y�JG ���iō�eyd�� x��t��|�$("+�96Pv���Mf�dkz)$2
$v��0��n8̜�eT��E�<�������k�{��t�|@-�hg̺���Y�'-J�2<��v"��8����2�f��!~�&UY���ߜte��<w�� ��h���gG ��9~���
ª�3���C�%�'���6���=�E?5&�U��=���Nw���t���=P!#3V���tҤP�2���	�J�%�<� D(�,G����!2u�U��IV�S�k�<�]R2����Ü!쥄�C��%x�t�𺽷����h?>$� zh~H��}��z+1��'�+��B��z�_�'�$�8z��1�H���S�0o���~
c��:u�"����ds��E�I=�*�+|?��F�~LbjAB1�����ޑ�6P�O�9
��y�.�T������M�t����hm-�7�E��1Z�3װ,�m��`ϸ=SH�v�ko��ɲD��V!�駐wM�F8 £�E��L���|=�m������8�,;�҄��g�a"�u����_pI�4��)p[B�*��z����'�s�F^-t�޿}^��~o��)}��O"����;�W�$��m��O������4E
���X��}q8���/�t�V��OH���h�/as��v�a?g�Yx$��>�X��)/yϯ��/�6�nIǨCDt��'��������O��������ǝ��Ǆ0�v�p��̃2����{zn��V�=�
��Y��f�M>b��9<E�rM���~�8j��n*"�}��]�ݷ���=��X|��d �������o�R�-�v��\݋����8Z{�B~1���*��ҋ!�L���%����8A�Ls��l}-{Υ����P��4*�0���G��[���ѡ/�;�^��\���8kg>f�6J��n�3c�D-M5q��V �j�10�)���#'@+H`&��l�w/mߞ#����F"Dݾ��n�O)hȱ���9�?bF�-�٢���k�qd����<A�W֑�wo�a��"Ԕ/�����㌿� ��Y�?l��q�|�d)Q(��2��8 ����ˊ��-?���qk=g��	/�I�x��BHe}�L�m8	�r�t��9�&�;J���r�py�����n�y�xE��b���`�r���Rp������61��S�$r*��=2����?����N<NA%��h��'t��e��l��`1���s�]n�J��w6F�m�#Ie\�i���
����Vj��Nv��P ���\���1���2k��1z�0aQ�ޝT@�����X�Y��p=!��9?��ٯ3$���6����͚��_���m������z9{���6Q�V�{wy�[H�j� ī��W�K�Ua�UhH���3��]�~���I#.xT%19	UkEa|
��t���C��A�m�&���B)�w4q�8��[I�F�['8�Z�����p2"�BQ���EB}!t˸g�d	���5�Kw�+���tϰcIʐ�4�A�z��kLy_\�Hn�j�&��'T;<�6�h{�گ��L��N$X��:n���u.�\
���cjFm�u�L�{�I B�/�_��;�L^
�{B\������
ό��*-wX7�
e,:����{�
�nSh�^࿺�����٣��ǁ�Y;�����֎�4�u�u�'��<��~HY�T��q�羟�K'ƽxW�4)x�j%������}rumg�����6���a��h��JS��M�R��$�w�Lw�L�/,�c����t�GT�"v��	T �9�}q ���N��GNˣg���m}�x��",������d$��s��a)��(qaG��/����:v?x#��:Z��C��o���W�?��qՔ�v~˰��C)�d��XMLW9ZB�#�%8�?���gH�S�A.�����M�3��Y��U�E�IY�CzMڔQ�@R���n3��)�si\nK�y1 �l�5�j6f�m�A�)���!��Ãl�/�ӛ�?G�%�Bꦎ[��Y��T��rPk�B8�!Z�=*b��<�������/��E� ��s��[k�|�
����V���?L��|iЫrD�kܞskm�2-;��zѓ�Tڂ���L�\M�
Ѡp��l�h�Ps������d��v`z95��� �8|�%R#�_O�a��J���PՋ	 w�O�g9ׇ��\�[��'4�������ִ�����u��"���i��$WW�ר��7�o����ZF�� =�ʌ��9��7>(��@����� p��E��3o�1��a�b�Î�7T?��N�<��h�k~B!��x7�-l$iƹ��H1����?I\ݮI�v�jp^����鯵^���N���6�]^��&�$�����;m�T=��3�w��g�q�;��A���wط�Z�I���[ֈ�y��0�	�i���6:\06��6*�T�D�eԹn�3�t<�Y��t�@Nz���Ю8�w��f��a|�Y�X�`Ꟊ�\�u��e����-��Na�n��_�,���A�"�b����ۏhG7�� ;!��qMF�k�v�6���QfzN�_���{�-�C�6����l�|LeU	_5z���!�[�����05&�V��[�$��/2P�f�K�ɳd<7���/�dj��}V={2^�y?ۮ�	���	�1Q�ܔ״��k2)H�����b�t�B��I���� �_��*Vn�f��c����C(H�!���d�cgE��e ��-������XT?��l)����i�7��yx��v��0�}�ҮW'�ׇ��<}-�7�a��|+�D%)a�,�͉��O����Yz�;
&���+�a�:� ��,fi�48ɰ)�vQ�Y�"��s�AK[��d���"/�]��豋�&@�Q�0��ǃ�\k�W�^Q��o�19)>D*a��f"��f�q?4��짾�Q�V�����r��ᐱ:g�A�eO�c�������������dc�G  �����{��k��5ZFJIL��=�V'�����W���-�!6�7��U�6��BΞ�����z���Ƣ�4���$�kF׹v��� ,S��.EA���E�3��U-�D��L~Ԍo�#W��U,\���G��ájm���'3��b�T��L��-?�"l����7q���A�%ռ���%�Ԝ����	�H��Y!P������̠Fp��M߹�}�xW��Ӛ`�0���jI�"`G؇�5��~��Z��6��eЕ�^�_姉6hMI�A�4w���~���ڪ�o�)ǻ�7]������;�������ֳ꧲]g��iO_'d:��~�ٰՀ�*>R����&A�[0����ϸ�~'��Jp�~Eo���&��b�|K�0���B55TS��ҡ���s�2�s���v�/��vN�QG�T��lh��ʩ�9�G��1�,g�a2r�S�nK�hY�9��C���xRHo��g?���0�b
gf�U�Vgy)a��$��d��8�u�M�\2?����=�?I��*�&}�;p�I1�mh.�G�<,SbJ&"����ZV�M�z�6�r�^��f���q�:�e{��c�Wy~Cz�I���L�A[\n�4�M)���V>o`xSy�@P�������|���)5.k._¥ŋ������*����_�ʘ��6*�E(����d��@튂�c��vK \q}<�w0t��!�p��{9���U���9�m7�/���|x��unaAu�؞O���)Z��O��-U�@�;���W9������#j\���*�f6:�b����QE�ſ;����(�'�h6����U ����}��t�ɂ��4,��x�S��dl�y��[���>¼�i'��z���{����*�s��i"2I%V��e��4K�W^��K�ʓ6�ǉD��c���Ԏk��E:���5�D���U�t�a	�m<�
xw�K�C}��0������{6ڀB�rO�8���9fzh�M�4 `T~��oaaI;*�"�EZ.|���s�Ibs�>�0���d�Q�l���潲�	�,+�g7�1ޝh��������' V���j������Qqͷ(�:���;w'@p	Np��:��;��;������w�z���^���Y�U�U���sΚk�\¸��.��b�!>��-HhGd�x��)t��]���L�*J��-sGp�[� .��$6������^��B���3����<u!�O�R��c�I��^��\]�y#�����!��C���	y����^W_>����I�%N�~��hkr�qn������6�x���9���С�-�?'���_���PD��D��C���{�Ӡ��-8��ڲ��{4���iQ�BC���]��0��tR���T[m,zl�m�]��׎�f�t4"}:��ކ��T�4��t,Y��B`�&��7Q���HQs}����5{l��:��u0�!� $:93`��=Vl��f���=o|bY�ZRPP߹�PQ2^:�������+�ᴏ���}�e��+L���/�zա�Jj�6�T�:������ld��##:+Z�^-����`K���VǕ�b�kj��kj��y}���4�ǘGM%?�`��2������p��	�v��(��ܮ^S��{,X9�e��SZG�K]uX��U�2�*&�L�'�Cp`�t��%k�����f�!��c���<fܐZ�6���R��e7rw�<0�� \���,ݯ�c%z1|�g�W��r�/��4�K���H̰�[��ʂ���Ћ�����
�1��N1��$�hX��͵I���T������)��Di8ڸ�2&�7J����cJ��R��M Vj47c�|>0W�	Wޫ�����q������ESH+��x_�u{Э/�O=��y�o6uݡ4s�j�]�NAcc��m�_)s�����y���b�"p@deeպ�������4["�!�ވ�,�&��g	B��ׁ����/�d^!�._d���B0���2���P{5�6��etd?L͓<������{6��~2\ʹ�i:�8%����9e�I��C5rT�򗬃ܑ�7!F�zb_��IO=E�jv&`����-?����3w���	ĺU�]�kQ#�b�e���_�!`Mi߾��)j�n�P r?�ş?G��ug�*��h����y�Q�_���f�EtV���H�~���7�S�k�<AŔ,>�U���҃y����1��=X�ᗦ��&$�$�>�m��A��W7?����tG;1�y�
=y�;:Z�m[Q1���W0��ѷ��@'��;���b���e)0B���#�d��>ޘOB�ϝpK�X˭ e(�]c�,g��FW�9���=HY�YPh��j8��Ѝhs���{?t�R!��HZR筡�9\�������?,�j��=�C�JG�J��2f��K:;3x��̞�|*�"�����:�wʀ��0f5& �˲�>��X��0ܷks�H�ؠgoDwn	ӆ�����[ւF����w�3e�����¨�mVU��FO��~:����^4)�R���}��XPT�d�_v?؊2��q�JQ7���X�׈����uY��)��8���y2�C.�a_���:���0_�b��h�?�²*$�t�H��8�tc����<�da�5�*�_(FRb��<�����Ȯ�|�u6��ǜ��������h=,���#F���L���X�i�(ݙ�F�1���0-d��0�ś"֦FFחn��-%:��*���4���onj.Dz�
O�F�έ��3�Ҧ��T����.D���y)��7C�3I��b���@
�<��.�j_E�.�
?�u��#&�W�4�p����-�1�ᵨ\}o+�7�"v����3G���|5�KOFf�_?�����w�'C�ksl+T��]���_��.�"듄��:����OI06)�<շ�a�c�_����-�D.ɰ5C�Ijؙ�AYS�ߧf�Y}h�7�Z��B�}�/����w�UL�mY����^�f�i�$������<E���^G�	`�g�����.�>D?��5y�a��,�Sw��oy�M!Ϯ,�M񥦢��3?+ʒ���l�4�|{gmڀ�S	����VI,X�L^D��+�;u�$TV\?���J[[����#��� ,3�;��um���z�p6_�Lj���n�b�J���t��N�$��QyU�8�f?�5�-X.�^[2�O�+��&��cW�}�f[�h,f?�t����t�%���Yj5QG�5pr�_>5O������X��� z ,6EG0���U# ��~pRXy�<x�C�Od�{[�v碲p�z��M��|��ΒO4�X����Xi���U�ߖ?	��_��� �R��O�,�x�ղM5,Հt?A�鼈������()l*t��l)��gRoӬ����/{��J�?ƅP�j���5��Qis��p5�&���z<��.��ǳi���v5�{aoѕ2v��4>�p��%(�t��j��.���c�E�s����$W߈p�,�!z)�|3�/�h!Wj�L{��CL����/��Ѷ��=�$�pȞ�!�M�ȗm�&��}�/����J9�XX����	�Kط��yOP�}�ؙ��@�6�k��p���"�y����>r�A�ݜG�k��hvK�X�!���o�2��c�C�s����,D�K�ד��d�;Qt 
����Z����T����p8��n��������OS�V5�a�#@�t�[�QX�����|����&�Sq��h�,h	���& �m4��e乷{���,(�q_.n �����"+���!�7�3k�<��?��L<y�=�###t5'.�I����ng�B�X��ʧ��]Oj]�ҍ��Nmh�~������Z_�V�")B��6��܏��؇�ŵ�b[l	p"6�J v��X�o *&t�_�P���}UJ�� Ґ��9�j��#x�W�ے�/�:5'�#���JB���V�~LK�۷�Nn�h�?E�Eݙڔ	B�09�q���������о��	ٟG���Ol̮�^��H�ִ���I�f=�d ��2@˩�"��6F{���H��l�6�R~u4u�<i���:�T�x�	�l/r����zF���\61L���^��&[����GBo'���gC�Jۢ}�>��b��ځz&�K����j��\l�8���'�l�k� �Rd�= �P=�	�f�I�a-j,��}��8Z��w>�0'��-꽀kܝ����W�p�g�S�cI�C[$�]�t��81+���53�6�<7�Ξ�)��D�>��<���1��ï�^Fn
�E��s�b�q��G/�-�0(�\��� ��Vw?�j��<F���ȗߦ��BLf+�S_|���|�^�楔�<�*�_\+�V{�0ՋXs} a�ܭ�Y7�k\�ڗ�{Cƣ�c0�4�%����)E�Mzv��y�v�Q�G�"������F��+d�i����F��	�x�fP��f62�[%PL���g�����e���n��_���ߵ9판��ͥ�U�y��͏�&Y�������G_���ؘ����{q�}�+,G�m\�6��6_�y�H��T�[���ꣳԕA�]�M�VN>aR�iĒΤ�����(���T���m���b��F����@�i��z��?���d�Bc��` 4e��R>:U�F_�!~+S������C؊���Ѳ��Ew���{��Y����/�O�_,�C��;`=z������i�.���6��:�:^�I�]��Z>����a�2�i��;�{m�����Vބ�N�����lV�>TX�ĸ�}�q�,�m��s�
�4�K����+�t_jz�5�k�Q��tm�Q�냯��-Xw��cm_p���Z�(��G�w���FI�y"����r;X���l1u��*�������V6��YO���蓿�կE�a1U�_�O�_^L~�
�(��Hc��K ��yY�"����q������~˫w�ל�H�}A	�Uݵ۹��������˜6������-��<aW���[ِ��w�#�_ؠ��\� ���B!�o&���u�����u+�zMR��T�|���9����'�~��zS���qj����Fޯ�����'|{M���wǂ��!x��~wD�+X��5C=K"Į�N����1j�4"��an�X�r���돳Y����M^Pg54�P]C��/<`7Gĩ3c�KW��_�K㑔�tâ]���I���cY%%ԯ��"b�)Ky�gIII�3�$!2I93����pP]�$���UUU����= ���(#�������i5��3<�n�Ą�_{�j"�ͯ]+$�:d��W��5H��r�������.�̃Wq��[p��\�5I��:3&��w���N9Q��4�6wQ/Y�2& ���+bY['s����v���*uPw%��P�P�����c{+��w����qy����M̼�h����g-��>Ӌ���ۖ�&A��\}u�m��n��a<��i���sߙ)X�m�A��q��n��*�Eh�o��s���>��*-)j~�"�OT���2:t������>�a�m�9�l0��ȇ`��ԑ��L�E({�\�D~�� �J���'���""U�s$�l�J~}����w���10Y=���H��JM@k��Y͎�a�z8�ȋ�ٿe6uF�Ǔ��s6�� ���sҏ6t��꠩[H����+_��#����A�����L�GGQ��˛do��ͥ�>�@Gֱ����⌿�p���1��믚, s��+O�n�k��Jr�=�}��G5�q�ױՖ���VN�$��i���_���0�h��cV���(��\<��dЈ����8@�xX^xZ	Ĕ���}h$Oz!����P|L`�
��&���4����M�Fch��gF%Obi�w+�&@�O���q
e�Ց��֑� ����#�Zɷ�`���~o�]�
v�#̢_��K�5d7���̢��4�������W�����Y(`f��������/��
��q]X�.���fu�uߺ���G��Ǚ\S����3B�r��a�����7��XE3���!�-�[Za7i�)�֤\w�7}T�,�Euj��b��|�=�
,hZ�uǄ�T�A�̔{��T��D3ظ�w3��!�;2i�ۄ�+m+0�y�ʣ�X�7ů���.�%Z��o�:|�/�쟷�X�Nߏ��Xe�S���[����Y��o4t�[:a��fLy؜d�h���T�'�N�s;�"�{?�a������ɳ�MR�#$8tg �7x
;��l[/sP^1u�7zBm���$���6�; o���f� ��f]��A��w�O� ��ؖɕo�@tN�w��޺�c�8���GL^����0�䮆pC����l^��	a���y�hji�$���wm��@)�r/�v��V��$5���EI5�Qk�c_'�� 6u+�}�إg�9��mg�"?)�BhH�o�50(��^�H/ڂް^&x����bS��^��%�O�����S}/�l]jv����'�suV����Z$�z��ͭ�^	�z��A��oE����5�$���j�����,��e��a̦�ݓ��le��X+�r�k&��G��*�7?	h�oU��d
=^5���<�^�ӜWC��Οtbi.�x��=�碬P]������t��
O�j�#�*�_N<�=u2�,�5"�I|1CBnËz�-V��[I~7k��B��B���H��5�oGPp5��婝���!��������(E��Wx��^�Bg��<l"������ۇ=����	P���\� ��Kd&լ���v�J�y���	�DX#v���/��S��P���֙�N��4�{P2�4J*n�W�P�Ft?
8�F��_]��ʂე,(��qP_() �i� ��;br�G/�2��i�x}��1^L�m��"ͤ�8>d�`���F)d���\�)��6ՠ� ��_(�K�D3�s�c�)�HeĒ�_"��϶�n�f9� z֢�U5�|�6�nK�C�L�t�Ry��!�X�)��Uggfq�ӢB}��s$ǣytQ���I����n��X�EU�!I�?M���W"a)Fi���t�P�8$R��E�
�P}W6�jo�E�pYۑ	~�J���=��eIn�Ja��<��¶�!N�~��*j1��~I��4���H�v�Q��5���}�>�w�v˓@�D��,�@JI�gփxvS&v�}Im!h\�Y�=�9��L/���3	w6{2$*����S�v���G>�'��a3���5�7�IQ�I2Y���=J��Q��%�}���޷B��*W>�v���crp�j��|���'w�!o?b��-r8�3qb�s�re����n��Ѝ���S���m��	ʆ� �I!� �+�E~�'����n�^}���]i��u��YYJ�3HJ�/	�ƒq�k�D1����
k%@v�L?^���ĀӬN��=���y�S�y��0/q��Y�1�����VGf����$F�hR�lP
`!.����v}��p{��P��I�7FgX.4�Q�L\.��0!>U���s���uv�Wg,�mJof)i�^9��T��c��9�/O �(Wb>H���ٟ�O㾧'��2���9�*|݄�ǉ�S����(��r��l���/���}����
Ct0��I �C�I�����Π�{��S�q� �q��c�F�� �Q�g�+�^��5�3�܂	>�c;����q��Hg��.5��aH�ບ|���TJ�l���ȼ�`"��l��fQ���ȌN�uz�;�Ni��Z�� �ݦ����۲7(��|��O\�o�Fs:�%%aU=h�t�������3��r�<h&{�#A!3�9�m�ޞ
|>���5T��JO� *w�w�A �p](0ZDĿ�x�!n�$
��S-]Mģ1Dd��^ ��ц�$:���iC�Z �e$��`$�r�ܬC���m�������v�4��f�~�l5�G�������ۑϴ��nz�wx�f����M�rl��\-����'lƿ$F�3fN8،U�b��Jd$����i�������\�7��Q1�c�	as�5��:b��x���AGhi_�ä�qzы���A�����A���0Am��=b^pF-�1TxC��ţN4]y�M^x�Tc�bԦl��>=H�{���L�˱�T����1��(��=���-ɺ�K�MCb����w�dyO�8a�k���H`c&o)�:��=pטF��:!�.��D��>'6t���y������~�?(��>�Q�����@މ��`q�O-����@2)Uȅ#�B��8�G�wO���-�wW�Β��M��ח���m�����+ܗ����FۺG!x%j�1	+>�nm�;�p��߿5�|k���Ή�[1%��G�?>���4E8���G��:1w3�y�^���[QQ�r�׸=ĉǉ2�)�G�#�Y<K��b�TDiL6c<.�T�� x��n�c7��ֱ��&U�v��0��
<,�~6f�h|�q�I�#�BT��9�X?s�F��/dp�2�4��&z��MԿF���E�W#*������ēÆ���k�I���҈o\1�T-�a}��ޗ4PY����!M�d<Гh�j�d��Æu����Ja�q�G����x>�#��@�M���I�P�u�����o�>IH��}^�g2�!~���n��Pj�3N��k[�]��L�Bd3Q�|k���_Xh�8���Z�����蜸-�Μ6��!�C��dK��A�q�pAq�q0B�N��� ���E��G)�:N�QZ��@��R�`	^��~�5���A�Jbe�o=e����K��c���,D���GqS��y/��	�J�q?�@>��_������f���2�J!{T��gC��-)O�L.)���Js��'πc:O�U���~	U�������S-�w��w�7��]����O���%��Z:���
�X�R�rӭcf&ދi\�4q����<�i�^#!k�=��a�$8i���E,,,��1t��Vl3M�P>Zh�9@�SԴ��h�8� g�YnL+m �v����q���^g��v�$<؎��Mr�V���9��T'D�/��E�e��Ɋ�Cn�h5n�����X;�k����M+mb��S�S���2ְ�%G�۪��/��ְ��"��Y��$�@:m>�K���ca���\���@���eE�7���ϩ�CM�}]���L452���z+�	��U�}1ʮ��s���d��@.(���]Ъ���GC����88G�� �pY�bC���4p6g�2�rR)qM7AE� !i��J��FbA��(�$����߆ʔ���֔�� i���RdP��p1W��Y(a�ZI�
z!�7���38�*�t(���4��Q{r:��W�_��Nom'�o�'�����*�/.&8�K��^7z*���F��T�?�^&�Wv3����z����Q{uJ�0θ�$�'壽���>�������g��xJ�%���VixCH}=��>O��'_���B��<���a0JL�=M�ѫR����w>��%=	�,��_�L�Tr8������:����[��N	�D��Ȕ���pQe.%l~K�)����!�ʉ	�A*��6e�irXp�����F���f�gД	��D��+�_ ~>�Q��/�+ٺ��(��i�K"��� l�G��JVn��M�:g�F�x�qd��F���5M���"�,�׈D��84�w�����l=�wZb?�k�c>��؂���%���>:�XZ��,��E���Ӱ^�V�̬ %\��-�J�������A�w����x�J�Ę����S�����Z�If��i;B*�g"��Z0�Ư;��)�����J�P�� 7iY������PL�=z�Y�K��ArA�ϭ�� ��ugOd!�60V��J�6��,GXǹ��{�~wT�1y�fְP�+��xPcR7C�=�������*�F�M+���Q[�t0�>��EZQA|$��j�(��S6l�D�9�sm����G9�в�},0`�AH���C=����י"466��9�y�Qg�g����
A%��4!�c�&Z�P4�� =���S�څ���H�� ��:�[�z1��a!���U3�o"m�������i-���Ǵ�Щ�8�ي��]x]� �4vz��K��bc�}�w%L���aU0 &�pE�}�##F��/g�'�Dpw\��96�a/���I��V�Z���^ڛ��!<⥝!]�?I3P�荂��/(yĘ��i7ڰ�0�D��ru�gzU�u� L|زbiGEV�
����8�v{�湠�%�@9*��]���n2M�k�R�E���T"-*@)&R� I��_�6�d/��GA17�kUi�3գ	%	�?DH��M�xti̼у��	f!�5Z�K�x$��ʱ��I�~@����j�d��\�� �*Z���/& ba�8�C8��9�����×��&2]��.S1�Fצv�vLnÈ·f���'$,�t����Us����B27�w�7�(F�0�~:!���>s�b}�-�����h;#�O�Q�|߶/�t@��<��_�4���1r���2�H��[�rءL�/����t��g��I��K��D��a�����kK6%�@)�",Gu赗l��p�H�H6;:���O����|fEٯ��`l��BȻwWQQ��'�ؤw������T=\jJ��������M7,?...�ރ��ALd$B�������$�|���i�#�dyY�!ҁ�]-?HÎ�b3򤫖8����Q�7*^���;��Ц�'��j�!2[R����B���GBj��hl-�=�8p�H=l��E�nIH���%8��Tێݴ��9i�O���Y���q6+�-���b
J4�����/��@��<�c'
��~Y�"��^���X��d(��Zo^�`�mIǜQ�^�*�X"Ggsư3�h�!�nQ��Q��1A����^y�nY���X��� d�.(����΢�m�ᙠ���fNхK7"��@�%]�?4���>��7�jY\gA�R	�h�{?�8dh�����%U?�w_��-[�EslM;[8��&�0��w#�`4����`�/z��ؗh���J�a��J���듧~�&���݋Ӯj1	q����(�E�0Q��bdM�B8��ِ�O�eSD�:#Dw�u�}�jr5(b%��~Ҷk$��Zչ�|��ε��	L�[��1�͠`�T�%�����(��
 ��v���/��Z��՝�h3�&^���L'�I�/��2��Jݑ��c9s_���i'�$]s����\�E��F|��v���#ۇ���� �ht��֚���71�nO�	}�¨yB�WȬ�:�;
zJ��Q�ic�$ݪ��������ָơ�a�VZӡ6�4��@�T:`2h5�
�!��g|'˺�\�_-�-�v��őU)�3����=����B�&�!R95��A9�8![IQ6W�lwH�ĩ@��_v_�z O�'T&+�K��T�r�_)��"�I<��aY `�R	ӆ�{����2��1����!��s�:�OE4��è��Y3����]�9o�y�� aX���*f~hQ��C���9��.�:t��4�_- �لi��z����Йn�j�g�C��x��vD#Z��������ۃ_ ञ k)q��ϣĉ�8�,ȥO��� ň^��]��u�Al̝��C�&i��\�+̳M�SSv��ϻ%�g���N˽��P�9l��]J>���>:W��0���d-��$�	g#��y Ђ�v%E�@=^O!�%NܫQ���s�]�ײY^�*�>�;Q&с���h2ܽ^����T�
�T�h�R~
��9ɱ�<���cЉ��h��I���$('x�H�ʔ��1�m1
-��hU�T��H��CN��pC�	��Hqw��2^���4��<��������ק�I�y ���
(S=���Q�Z�P�_f��z�Qf�B���d�rG4��y�4�	�(�@�R�l���	 ��5��#�k�òD<�|pC0!�w�l��ys%!TQ߲5�� ��_?���H�,��OՁ�RL�x�J�M����ס;z��������4H �����C��	�}SrZ��v��J���:D*�lR#�rV�C�~}�s����5�����2Y�`�E>0vxS������ꊳ
�+k�C���$���O�@��}�g;60g><9�pހ5�j�G����������L�ң�P�������>�y䭹Q>�P�`�N..X�v��GZ�ˏ�oP�����I�̄�mk)�X!%:P�9*a _Ͷ����` ϻ?�>_x܎b��g>1#�~8�������:*NpgFn�~klz%�����D�Z�]������yE-��ߣىn�҃�Gd�#?:Z��b䱆�i�Y�!Q���<?D\5a�kN<�9:��[�ϵ�`�x�ni323g��z{E���d�"�����>1--ӭ�Zz��M�4�`1p�U����Ǭe����Qm�w����Q�㤢���ެ����O�/R6	 ��{zb� ��A�N���E�x8jj�͇t$Ї,u�;
�ɟ;�d'G��1���-��\�,`��(��w�a ����=���劳lz�@%�;�?0���[g��?z9濧���r��3�MGjuJ'Cl0�F�pk�HIL���#�b��~9G~���b�N�� 6����7��kL�#�+Q�j���������g�TGd#,�ؼx���k1���R(��V��b8�a[�W�Cn �ߗ�5�ڧ_۶S{U���Q���Pn`q���1��A�8����|q�)O�>�*�*�e�1NC������5�y������[���󮨏 Q���N�9���$��wy`xgɅ�6�p�k.��|&}������ 'gR ^����a$-Oѱ�wPl����i��d��12`h�̆�����uf�@$� Pg<�1�{����G��ї1��vA�o�L�2��}���,��Cjd�F�`)�4�z�/=���n"\qN�{��^�@��qz�5=T��ܞ�"�	=C�'�/���7S(�W5��1��z!h��8 �Sn��F8� F��_4j��k�J��C���h�G�6�X.���`��v��R`g��](Q�L\M�fW@6�[��َ�_��_ƫPyߛ����@����%�b�����G
�{����î������o��KO�	�qP����?�?�;�*xޗs)P!��@�7��#�%'��#��ǁ��8H���"�:�t�[�jX�d�˝(��DT�T�c���49�X�T�08�̊Fb :_o�K�l�`:,_�n +ͺ�P�m� ͠c��y�5�VY��0P"�/���� ����,�<M���������-)<�F�E�Z�d3���!�(n�+K��/�b��֯3�?�q��Z*�n=� ���'Q�{��#�р��7QFw�3����h�����s����ȃ��C(4͢I�~x�k�vT@����A�U�W%Jͱd�6�l'`Էn�\�E?����φ��|�p1����ɩU³6{	�EO��gm��r���T 1�Z�z��pP�6���-�2@i!Wi)���������T#���I��h����K��ö�چ|�X��i�Z�@VЕIY�#���qW]:Qﴨ��p�ݘ�JX�����}�; 8� ���@Z3?U��A�	ĂU�-d�*���-�l.�N��C��t�dkX�:�2(�4u��VG�BA
�75�GH�Ϝh����1�*�x��rNP��H�6X��BK_mo�r�A)B��hsi68O({1�>�;�-�d7.x�������l>��g����|��vT�yL:��7�H1S�D����e��K��������(�2�V�@�� %��� /(s	�@�!t�A4V=H�a}��0J��t�o��L��6s`:�ӄ�U�ɍ7��ЃH���yه�ݹ�xH.CI������v0�
A�D!��Ep0��Hm>|d�C��S�w����J�0��a�F$�3A�=�1��<LZ)ش�q���0����\W~"~�b�g���������nTf�\��Gg5Q
$�^��|t���E����A���Ľ��0���*���UK����ߎ	=�����1vnr�J��A=�j�=�x�-�s���������Y�CU˂G�^���y���\�t�V��U\͌	mc�B�#��uZ���.��~�L7Mxl(Q����O�DjA(Hަ<�/�[H}ʕi��a����Κ��R{�k'H���&���@X�T6�}�1�@�n�O8iÌp���O�x�5�c��'�ߋ16���i�ؤl��Ζ;%�2�]�<h�I��D���A�ɘ�}��Gʇ-������N�@9G�f��j���g2%#�NDj���!�s\��h�ꡜyJY!%��E^^�,WpdI��))�j�m��m�/�o�0>lz`Z�n�NLR�J�"�{�ƌ8�H8y�F���µ�dP._Z-
>������E��a2B�����;+�^�h(��S7���A�ؠ4�>�W�'�x4��`� �B?��N-NG"�n�7O��f��j�K���!0꟭�)�A���m�\4d�uh�;#�D)���~*A-��Nh��`�ڛ��1�ü
���ƿ�=j�Y��#�,�3�W�X�*1��@i�r�I&�) ����u#a*sB�����B��	�ʪ5f�5TE�ں2	n`t�����U���?u���Z?�n�@�T"L�Dٞ�y�h�`;�7�V�ӡq�L��bI�ٟ%�O��aч�e����L��AГRo�8�;'�9(�sz�<���O��o{��Ո�*ߖ�Y�sM=�#����~H��	ؠɈ�7��>�z�ڂ���aL{ke3��TJI��?�ݽ���"=T�T}q�Q����HĪG���O�LT_*�Q��1.����%�ק�f�����j_�F�`$��S���89кd�mlao��_�J�0u4���/�h�1c����������e-����܄�t��׹�~>͵�Qw�C5߭HH�vh�|˧sE����IW+�ި�
���?��������p���d��i���G��c��Di~�zԵ�C���9�,D�Ŗ�b���IT�x}y�.|Ȓ�
N��x Q�)Y�9)�S��#���j*����o��������Js �$�珍tΪ���7��ef*֖�X�vnE�qy���R�?.Qf��~G ���)w��,y�`g�m�ʣ����D��_�A�(KqK2g��v�}�7�M��V�u��=���}��}������S	8�V�0����E4%9掉�=�01�D��ꯦ��ᄘ��>�(���D�)��g������[O͞�瓯ܩ�&�YUL�(�a��]��m��z���.�ӟĭ�^�w�Q'�I�1h@�q�J�B۫WG��0��f�IpQX��/���@O�7�����]�प�]�׎�Yyo`%�@⤑�D�%h��e��d#����̊K�	�l�R�����q���8����Z��inƃD��9�3�Z��p����$����Y=�A!�-��H!N<v�v�T�;.��:��8͌I�I��%��H)��[������m�좊�F�����Z����phګ�-C�y���u=nb%�:��8U�Կu��1K�"� �M�y+|/�`�������u ��/r<26hJQ$���w�h�W�F�C1��F"���
�4Q6������o�l��	�J�;{W0ɠZ4��'�#�[�`� ��~Ӏ�����&ڳ��[�I��(Pw�u\U[�i�7رB�ۓB����x�y��D|��8q#[�*/�7��b��m,�>��*�!��t� 0B�M#7&êe���������[]y���K��?��e���{������}=�8s�MM$�p='�y8�נG����HS�{H�;m*:	u�ݠq�ø����u<��q���O�y<v��"0�ơ��@$���m[,��LͱJF#��5���Q@jsFFL���DaJ�/+�̦1��<����%��Do=�:���1J��HRW5�����.۷��,�(LBF�V"։�?]�"P����D�vm�m[+F����:I�{-̼�ri�c��������;j��6j� ���1���� P�̑�M��a'`�LE og��6�
͡�����dB�>v�2H=M��Z�44C��8 r$�ӆ�pn�I�1�i;LT��^R������ج�T��Yn�-xD�v�B��l�L2S���@�-�Q-��� ��*�B�PG� ���Q�1"�L�a�g�0RǷU��*���G��N�\i��T#J�Ћ�U�׼�d�-7�@0��'L1$ףA�xfy;Q���]��S������ŉ�=�`�h�������a�����Q�,��B��j��c��1�*GEe����ϥ�ɗ�	H�҃�s�Bh-]=�X�}�����^��/Z���=:ŉ�"H>��l�x�\>���y,�<ϴ>:�˾��%��$�d�(��>��ݭ�ev��{!�o��R�4z��6��x���a�d��OH*��:�V���,e��+U�r)�ؓ��`ޙ�����IW�g��qDo�RL5���P�ޯ'��`�6]h`��7��~���{��>t�=���A#p��w.�x��o�i�@{&�����A�=�RC"~�R������ `�O~(6<�#D\�5�]����R��y_g"
D.��BX�I��%��U�<��j@<��Tڴ,X���$�a�p��X�	3C���\<��Ru�r�mi� �uU4/8��p1��<nwdMHSW~>������TOU�g�}��t�'���:�]��d+�H6����W�4�(���EE���@#C�ɴ�"�f(X��&��9��`Vk*�V�߉F/�wf���p=�����~�&�@	ؠe�'T�2$���Y����y7�z\t��-о�B25u������A���ag}#�ѳs��|��������'c<���(ly�[I;Z�6��
�G����^�0�	��M8O6�]G1XԠ=�ϣ�b���Qt�B��}��6�PHZ��q�*y�y�qw����D��F�Au~
�/��S{���B\&�X��J��7��Y�[���|�B����m�~G�$L݁*�m~�78��X]Db#3'lG�V�`<R��X��շ���A߬l����J���&��V��l�In�t���jmRT4�2�Q[b�v���{WD�5�d<�� [�6�g�4��L ������%�ǭmq`�z.2�H }4�Tt8�Ѵ!O�8pB#%��i�q�ĸ�S!ڎp�g!h�A�#�<���g��ڪ��@Jt�!.;@�!ZZ%�C�5b�If~O��U��5����vg���骢��-�@�ww��C�������]w��۠��-�Cpw�÷��2OӧKvU�}��j2V�"��=V�#��H����8�e�I�A��x`�,�}�'�k̕J���#�=�J� ]�N��
�}VWu�`� 3������bm� ~>P"8�+�S�L����kK�:H�^���B�2�{3x�bB���ZG��e�.�l��D��M�`��1��b�h,�G�˒G�5���f����7d��'�{��xlT�u��� �Qg9�U�*ÿ��}��mϪk��Q�l�I�-�r�"*�8\E�)�C}��K�ɸp0Q*�������g�C�e�g�,Q������}n�i�A�����*����'H�d��Z�#�O~/�����&ΚW�")iG����YJ�h�9e)2���>R��hD�#��G.��T$�)lx ������φ�9bΚ\�\��H�e�%*�a�bm(�Y��
Ur��tr��F�@���*��ߨ!S2�(���usd���y $X��"b'n��C���Vy�VZ����~+��D�!E= �r�n�0�Y���1�0.Ґ0͟�S��i�D|�6����j��U�H�I⛜�X�۝C��r�DʍG�/w��e%\�t"i��!�j4�ؕ��@
��t�3%���p��w��\_���
�{�%!>�˥K'U|?||,��><0��ߢ�P(s4�(	WT���b����F���y�{��Afw�}��`�c<�I�l����^,�CRh�3��M�4�
�a��e')�.�Z s���:�*�W����W���s��I�����Xt3袝~�B�K$N�EnڱBwOOK�T4١�wc_ɖ���8���jA��]Am�ܓ',��|,���Ƚli�=���J,,�͝_y��ca-̫JY:��#d����;���M�7I�s�k��c��ԡ���/��JݔA#��
�[��/���������?S��Q�`oZU�_t�S�Wyu��6_]H 4\���nH�)+�܅A#z��!4�H�j.��E��(;���.`��=V:u~�DҔm��O�#;1ռ}Z�{Z���/���N�53\��7\�/_�*`H��!�o�"�*jK�Ա��w�Ů�B}#�x�ȩ��Ǚ��]H.����g<�Rڙ���1�+AzāI5���1n�4a��~V����M~}�Q0F��O�쫞�oױؒJQ�*�i�p�UiH*�2d1V�{��b�X�.t�5^.�Oݸ e'-e�/G{.����������p*Ѹ-f�Z�EItx��J�tH~���Z6A�0j	��6��@�7�).'Ky\f\cd�Jg��c@\L���y9��>�������E���X#�SG�V����7n�B`���8��w�Σ��.m\�U���a���ɇ�#������O�Qn�G��j��=��l^#V߅�D;���4����i3�W�W�/h�5�͌��Ӽ�/�|�-�uu���\�%��l������4 �M4-'�ݥ;W�DKG~�?�Z'>���U;�P<c�A8��1�#ϕ?�3���c�����>��E*Q!�'�4����FXǏ� ��=�w�M5`22
�p��f��9.�j��Sx5QQ/����҃(y�0J3����̀��UA����ao|8�M�?��]B���z∻ֹ/�?�"}nye�� ���h����|�ʀG?k쇋M?r��	�uz��/���x��a�ˎ\�E8˵���2z�n�u�ď�#T��~���Ŧ�z�&�`e�� ���[�T ❯&�ü'ɴc(E��'���@s��I��f�E6���c�ǁ� ]�s����I�ַ��2�:(�4�,�#�`�"�mtlDK�д3���\9F���wC��e��z�K�dϐb�WQ�h�v��-o�v.�L�*�]���%|_�I��,7!z��W	�G.�v�Jm?���u�D���SQ��оj����S92NV0t�0����-h���������s:ؿB���tpɟ�`@�S��`��dܳ'eq���$���nq����fB)��)ZO�<l���-�HЭ��s�5��z"M��#���|��M����q�7��&u�c{���<p��h�^�*��kD^�q���3�ףE�����{�����|JW�}�9�p���ԝ��,�5�g�>��w.�z�W���뷔姥VZ���ϫ(5������(���$�g�׼1�^6��65E�vޯ�#��O7Z4��f>��5�������-)'n��ފ;�ǯdC�&�[	��ڹ|a�{H����x3Q���Q���@E�g򮪀n��T#����BT e�[�V�~k���]P����+`\���ک��SٵGC)R%["�V믶�tj}��"�#k{�wd7���I������A"Ӡ���P��}��ɴ������DV�
�˟�9�og������M��+��s�D�LK��|n=lafՖ��Z�L#d�ڷ�w����[|\x���O0��{�_
��%7�#�O%yJ���~jɧ�fo\���6���(Z}��bwSF��]�p�{�t1�����vi�b	4"�֫�Z�ξ��"�L7j믌P�1��v�� ����N�L�R'�
T L扩(�L��^�O�k����9G�ڴjm��ƈWX>��@~��L����\h�:�:fHW (�ʹY?F���6:�{�E�}Q������tq��Frrl)��i��}�.W�8n�Ahnqޟ��ΚDVl+m��M�F˰���U��ة�R����U�������#(h�%�v�V�B�oîE9%v����u�O�"!�-l��$���+�s��DT�~.
<	ñ���c%�p��17�������hvG����5�u�aR4��v�b�;�Y7�y���ύ���%&Lh�
ڦ�|�K��P*�f��n���V�qvlz�z<��2������a�� 6�|�}��J�d�N��^b��2�
Ӽj��;��K ��y���m<.<j�8F�N��Z��_�
��E���ߛ��[�G��)\�K�#�e��b�×�����vM,�v��_���v�0�ԯ�����M�U�j?#�VɆB]�-T�
��{i�.�b�x疲//��~k���aB\bV��Ф�w��ƶ��v.��~<5VO���g����*M8mH�8��q���u��g�Yu��<�i����7"J:���T�����5>���������>̒-��E�� [�o�~��i�!���)��z�豺�g��)G��S��'���No��G���4�5��0��p5��f��m]��@��X��i)m�l�Α�a������a{�޶a7�����U����L���./�\%�}��A��������B��x�mn��!�H^Ʋt�v����2�Atlu:�>MRY.��O�c� c�����l)�(�k�3򱶔�����F�DR�������$9^1] 8'��ҡ������ ݢ|/��p6����>�q�B�mк�����E��s��a�0{Fi�˩���q���dNֵj�΋Y7�_%��;��~�a1�t�,�E�`���2L��z���[[��u]{��V�˨�Oǂ�@�i.鋋)�ٙ*eAc���1������	�t����߮�-��?�U9U
�����;�L�I`��^DkR�ԯӦ�zAM��}�A�ޯ�������5cv��	@)�%�WwX>�e�)���F�\}�O�G�i�U�m�n	�Y����y?��v��'���X�+��8\wm��\6V�T��f�#��Q�g���� �\c�/	�Gs�
r	�/��ܚ{?�ef�F)jk�Z#�vfZ4e�ֿ������+�l�K|f�<��)&z]����k_x�8v��0;S�.�l`P��߇�I�#,����U�;p2�����P[�oe3���" (�`�3����W�,ﺧ�/�������K[�X�fE�F2�_��d��oR+��X����)���P��+J{�G�x�TH�r
"'Z�8��?IQ"8h��$L�����pj���[�!�v��s����a����H*�
{F��}`pJ!πi�z����C��V�UO����@���.WҐ\�1>���/!��7����Ӑ($ŲW��e����·E/����6�?�*���ٔpVlX�8e�B"k	 ֵ��W�c��qq��ĸ\ya��qVv`a6�ނ?�(����ڔ�~��r��ia/j�&�t��W����+~�(9�	"�*{��iү��~�6/^����������T������kd��1���m!o�MqJ�Q��V'�QP������}�u�
��k�}�ڜ"[+1�V�;B$<5Yɓ�X�Ή�y��h}��oRUc^�V�d����,]1�ӧ�ʩd��X��Ҩ�J=Q��5��~��~�W�;��=)�Z�QvP�{`�{qM�/6'�$�M���9o�)	,3P���*��1��-瑱TYh���>"�b+�3�X�6���*u�E�O��L%̧�$��b�#��x}���ܜ�hĨ. 8ǲ�U쫕�EV�_>�:U�|�ѾD` ���m) �S�j�Y��91�hP3�Z�ς�p}�]s}J�a�Z^�����
ݺ���ւ��Bܓ�#�63N�Ӷֱ-l������+��MM�3y����+7��b�`=0������1��X3l?����,���)-�4FR�"jQ�#��7��O��6�]���'*ѧ���nO���kVu����`4B��=�/j-1�|��~qA,��Y����O�L�1�����U�������z����E���ö���  $ ??F�X��]:"lj#_� N���G�*3_{1�/7�u��e*"�3#^�qV	Hh�;F��Q�T�t��KIJs91�	�3/�W��&��pG��RMw}�O���Ǌ��w<��CV�Y�E~�| L���寠��3���*wG�U��z0A��e�7�kE3��K�O��	-N6����;�aT�d��.�������%D��k@���9��YhJTqR̎9x$����L�ؤ�z C�|Ǉo�)��G��YX|�#G� @�Si
���W�!��!�n΢~�Ӛ����>��uaY�پ6u�J4X$�7�JO5̥�����{��L0IDȓT���7��@�@����WJ�)ȶ�$�[�����:�	��h�.���!�mPcY�yz^�����*�`�6�5��^�j�]ø֓4��W�[�Vn^)DUL�O��2xLa�]��_M0�Ԫc�;����p�)$`�P!VH�
ƴ%�P!�:��%�v��?bLf���
�p ��=z�2���H��s
t�<4��vK��̪]��zC��늢�ݝ�iJ��1s��M굷6_��b��I��
�x��1����h�B-ub5�m�}��A�x��Ո��z(�����Ŭ��!�\�-Vv@�וm��)y�WP��?��1�^m��a�㺃m�GyV��A����y��>|1CV��ލ��q������ꦚ�.�H���Zd��]%�q������#8;�TD����"2 ̫��������1�����!�j�ypa��n�t�;�=�_D��	m-.����}x�}�v�'�
2I`�<���P�`�f�V�^T���Ev��=Z?��P�b�>F�@1�N�JV�WW�ZL���� ͘�(Ò�)�E��v�B(�<�o+N��Ra�>U�M�q�'��Ƶ,z@M�-C���`#�e�/�~*_=�C3a_i�;%t�XY�OMI�Ŷ{_e��'�=rN�[��P0G{YE�ze��:Ѝ��u|�?:x&�063K���6��*����,g���C��̅`�\P���K.�f;���k�e�,%ު5�M�c�ۮ��i�![�[���S�)�����F�фX�Uw[�޺���/�q������!j��atZ(T�����ĉ����H=\R�Zn�o��H��O=*՝v�,�XiE���.F����w�E�1�(N��[��o�L�wb�1��=6����u��4���-Vg�Gб] 0���M��r|��x�%�H�9��&�Ց'&��ç�^b�*r�q��m���͂;��y�'[j-]`%A�5GEv�ը/u����n��7�1�vU��R�I�?����Ve�{/��!8��ZE�o�~�]��&���_������&��w�JL��!=k�J9�N��8���q��Ry�׋aT0+�Q�6>��gj�;ץ���:@�k�K�A�k!-���x�,��z�����YD����(#ծ��,�z�E�p�|�e�$zL�Z5��
*�,D��Y���sv���DF*�f�~r'*��Y.6'f�Ô~���E;�J'� ��H�Zō�-Pa|�q�L�eU+MAm��s�V��|��i�y1m=����jʸ��;!hss�$q�&5N\W�jqs�~�W��q,�3�����-���� �[���Mx:��Ӿ�����ùyj�M�_c�9�ϳ'����+P�sO��^�T�)|��XMlp t&�B�:U���P��L�vvb ��P�������A��j�m\�W�.̷�]�1T��iE/TMD�|��z�����"Ie�(,a��\�[��BU��1�����0��S�}uߨp@����s ����7pC91���Lcʨ����ԨPd�jF���>:��Q?�ϟt��F����� M�Y�O��5>�c�9���醬HH��t[9&Z�(�&Hd�z���|�>��m�Gh��ԙ�A�U�(���u$�(��|0ȯ��\u�Y���ȹ��=���_��'�hem���&��;���*m9c�b�}w��ک�������s�U!��!ݹ�^Y�{��.�V��٫���f`=����1vkˤ������&xi���'���́0\)I8r�`:�7���_���;A��"%y��c�u*|����I|a~�Q��i�c�q[,��wZ�+�*�3��9w�׀k⎇�`��6��	G
Z��C�%��8����W��ř�x2%��5ʀL`�}�������|4H�=�9��H�X.�L6X*3��M&)L���L�	��T!�f�>~�j���줻!����F���C�:)�Z�B9����/�SW�w��6y����x�MMB��� (H�H�7�w&�BH����|~�
UE1��+V�'[u~Sr�h��6��JJr�V�&���a��ɜ�wg�6�oi�,���79��]w�B+��	�q� ?�bH�T�������*�0j
�	���i2�!�WK�J\'�>?��J�,c�oW�Z�����j��!%�����a�'���a��"8.�Bm�>��� =� =�gJ�!��,3�Oz?MN�����;5;<X��v�y�M�N���"g�O^�;ZvR��]���Xڴ���x���^	C`(��	N�������$F��.����)���6�C��DR�?HP���lN ��o>�E���s�|%�?����>����U_��Y%v��s��$S�k$�(�g��K@��U�p
��c�:s�/z��~�Iy#~0Y�="h�"���A�x�>Q��a�΄����^$W.��щ�(�gv���C�Aj����̷#�z�Y7�ꔑ���#6��ۆ!%>XMk�/S)pCg�-e���F��ˣ.�+�,�yD�+�(�@1���@���{���g�Uwz�{��t�3��6)	�@9�'D
d�Se8��{��%(O�%�H ��}��;�( �l���qy��3��U�S��v�ڭ��۳���}q��y?�I:3~sye.�s�����0]aFb�ϕ���f�#J)�Q��$����F�%�v�^vb�5����z����73�j:8I��D?�tP+�?ē�z0(U�-�g����RP�X��O�Ɗ�8�ۆ�W���קs B���QS+_Zο�:��Zd53��W�t�<��Q��~��j�����<>pF�U^��n��cR�Kn�)�џ����q�M�֨�+uٟ���rςy��0���6�Y"Zo,��� ��q&xp�un��c�oiS�a}L
z�ٶu��c��&�����W�1Q9t �}�,b9n��Q�?%�<�88#�� ����F,�b|$%-�.U��!8s��Ğ0v��E�Ԑ�x��ErMZ�D�ET��!5f��؋��^a�kzE��'�PPɦA�#K�]���r�Q�׋�f���B2l4eЯ�g�N��*��.EDD1@-ɦ�_���?m����jKd�5�I���f��B�7
���lH�}���O���<]���㔧�[��}\��Ӝ�߾�j�E	�+��*��J�#q���ϣ"%�(܋`��n]�]Q/(E�/dV�����0����&+��b��$8OD͍��ZK|����� w�J�@H��B����%T�>���-P�:�ä�'��2h�D}ɺ���Ͱm��o.����\wE_��W�(�'�-W,���k�����t* �,8�3��B�����Ğ���ճw�I����[��jR�ea�:5���d	]��
���iM�4��]F�23�jP��i�z3C2�|�K�� �+Ţ�+�髋��W�ĺF/��\'�8H��0<6��x��Yqee~raCp��N�I'�AC!��S,1���T��$�%D����4�?��N.a���Y�:;­�֮���G�c�40�)o#��J�(1,�^F߉��X�-a�B��F��F��� Ճ?����b~�Oo��{�HY��W��~/"2N��z{�Hk}"W��)8s̥�bt[_�z��$ ZɊ�H,g��k��u�N���@�-@ToGA�U!�Z���9ƛœj� �=��EF��o����B���\E�A�����E�ϟg�j��p'#���������,Z�O�c��y�$�J4�ƌ��-ė���b�Sd>�gf||�Ep忷6�AT7�%���a�<� ��D]S�k|n�ub�.V��;��DD��K��ݦ�.�i|_�e���q!y�&Jtf���-6&_^�8F�tK�i��5g7�jk�R�}4��OO�/9�?�{a���~Y��a~|�s��&��	�s��K���b�'Z��΂(J?'?�y��k9�Q	%Yq�6���OU]X��9�c+*]݂G�k��*�S�>A$�� ���Y�D�B�{��[x�a^}����a1���nQ޺��=�{w�q%Y2�U�⇫�%�����aΤO�!lG1Y;1������s�Ǽ8¸Š�S=Q�>0��=lx�J�?��L�4$A�wz`i1 Wp�����U���,?�������g��o=eHL5�k�3����_,�~�GE69Z�StG��,���ڨ������(���]�BL�3��U�P7�b�z���hrR��sɆE��Xӏ���.�7�L��Υ�Q鄤���%�`{㺨2�"����?p[� �y�l�VmL��
��P�!r<F6lr�q��w��?YC
DXýϙ��N�B[d���������) a��_�[��P���4��)Id�h���ZU<�MF���?A��#�;=���KsD���O�TF�����&!y�������|y�� �&�����k��M���U�`v=Ѩ��thY)�N_U>x �I�N�0���G��z�D�5��8)Y���,z�ؒ���>��C����ꊄT7��eh�3n�EP�h��F����k�2KZ������+n����Ǣ��*0S��V �{MBhb�#�4��e��AJ���&��Ϡ헂�~��{�P���e�b�!b鍹������#TE"�aha�,�N�,?�#���iL3Fy�z�}gf�����:%Y]i�U|e(	R�c�e�O�r4���/҃~iI��'��ϊy$��u��)���5233��5���4Y|EɃ�e����B��S�զ�@�7i��8N$�à$�R�<M�΅�B�2��"�B��R�d�������r|ٌ)���EQ@��7��/:�F"YtC�����A�Ý��ɛ �Y��n���?�`��)-�%k�j�c�g��q���"�q�+��E}(��<vw{���TT^� nҠF#̶���Mx�V5s�o�nG��D:Ku|Pq�����}&	��!�p 0}Eol�e�<�r�T��~�8��\�UB�MP'��M!Ã�_�ʖ<b���d�����|�P���'��=�S�I��U��Ex�d+Y�=WS���gn���K1�T�\|�f��r��i��~�F�U8�tD����>�#w�	$�����O]�h6G
��M.,�1������ԛ�Րp�U��T��O$���C��|Y�������D���t:�َ��P�>���Hw�$�!&�n"D���c���aq��'����4+��6�s$/e�	�ފ. ���ߧ����K������ϧc�q�"��Q%0�� :���m�;Jt4�o�.��(o�����ηtF�g* ���Y�<cɬ��Ter�qVeX�(b�� E\Z�a��H�ArC#���lyC8�8^B�W�(�Ft	7���Y^�#�j�Tٓ�8ZQ���l�u��紤2`�g�p���0n�̒��ȤAG܎�e�g�K»�^�Dޣ�����$�6I��r��={��#�>�	N[��d������
�AB�@�Vlݷ��,⃀� ��(�O�9K�W�10��� ���F3�����N�?0�Ga\�������r��^߼�dkK/O~��(��w"H��I�"��N<�8��)�L�﯇�&�{������I*Ĉ��tث���n�A�#��K�[��0�w������5ڛ7p��dXS�K��Hƌ>"K��^ �b"{^F�"잾>x�@}c
�"v.�e��~���T3�޴��&zx)�ט�N��zH����F�Pc��Z��� ���׵ɏi�j��Qs3��+��Q��`������U
����n�5�������)9�!���>Hw-��`Ez0���X�%�\�Ņe���3X��6:����Y�9�հ3�����ƚ�6R���O`��&���;�u}��,5<*���YqQ��<e1�r0�w<͚U�=~���*2�#S�P�s��j�� ��X/�����륎bw3�%�{\bؔ��'���9�T��\����(�no(���,�'� ��I$+�ݼS�[����Y,(,��_��V��1v�+��Z�5j���k�`�*�K}6�P�4�&(#�d|	����(^�'�`�R��`!?��{��|�lz�4���e�����_olw(���Ȕ��5�bQ;���7���£�)����^�J	��ݢ�f-��֢*����]�Ai���n��IG�bDH)d��	���T+���3BE�0����ɨ?�{���R�s�"��x��O��O�oM�'�#��Q��r3F��0"��
�)ѕ3�T!�	�r��|l���3q��i&�^��C���2F�}�e"MO;㒸��}#9N�j��ʞ���Ƈ��J�{���ty����
���#9�C��c�G��VWyn�׬d��$V������18��)֙X�u�1��m�c��;H�,�����Q��"=��QF2ذG ���]n��[Q8�i����(�U�ƃ�� r.J�6��J:��G�� ��}ӱ�h){���b�j�:׹_X[>�!Q���=�_rlÙ�4��pW9՚M:�7@I#p���ɑ�ظ��xb������QF�m���m_�Yc��~�#>p)���XxO�#�c@$	�l<��o*��7Lx���	o�666�K%#���r�q ���i��o��rһ-�}����#H�|�A�Srr$esiY��c�{LYN�$�rW�{�aB%3<�ٗQQ�����@�'JɳT�����lN��u�퀶ds6��}/a�>q^s�z�$%�46��Q���}�b#Sg�]��Q��@l	b�������շr�T_�ݏ�X�&0��ˊ�=|)}���n���,΅kpDs�Bi)�y�$0
v��jb;t4Ѥ�iѭb���
bOJ]��x�7iq��b�3�I�ϊWڜ�^��s��Xv��sD��ŕ<_iq��T��2H�h�MH�YF+����H'G3P[��G?x��=��|��d�P����h	�ʋS�#��,��o5��]$���z�}i�s0�
���9�������}�\�������n]�R?����!&Tm6geý�F��UN��1�i���q���,J	z����i�{�K�)��[S�
�28a(�fg����L�p¨e�Fdݧ�_���/b����]�z+��➘c�,{N6'�u���g{���s'w�1^k�W��1��Ѷ��F�.�2�q^`c�7��`��ϤPW��ɷL����(yx$;U��NX>�>}�'2�!�#áрXik�&b�l�K>����C��xF��)f�:����B�α^ñ\3�n?AG��נ*�x>p�@*W�T�6Xr��`MA�_�hq|�/x�~���50Ǻ��!�oըX�6n�p!�Dn�M���,�{Vp�2�]k�FL�a66�L�V�4�OX&a[��m���)�bP��fę�n��Rb��$}�h�h㺱q�= ���p��� WY�"�����(���Ս���z_/�g��П�!�9 �,N�+�^�;T�*Ryx�򱿰����Q�4ָ{�,qG��D�"�O�+X�#q�p��a	]5����_��#Y��j�ڣxV~4h䌦_
�վ#]��.�%�zv�Ӳ�m#ʊS�ز~-cF���Ȓ7Is_-.R;д'^
Pb� q7(B�-O�TժO�^�f$f[i4p���3��?������S�3˺<�Qcpy���2h�fbW,己:�a�.H���C8��^�������mR���a�g��[�s��4B��m����UC>�8:�=�*(\�ͬ��mn��fވ�G ������A���:S�I3,_"c��,�&hDR���v`��f�oJ^G� �
�lt���3����u����3�>Sm��Z�f�k}5m��u<P�w;N�� �DhV�t���M�c���2��q>@T>�Ss�t�_feF!��ő�j��Q�MK�Ul�/�36���;\�Sn����U�7=	hf� �q���N�B_ue�^����]�m�kVGWr��c~if,�=�UϽLS7G�T������}o�[\���j���F%i~�
7��|�ӡ#嫇�u� ��?�*T����\Ung�O��no9n��SO�&��8�X�����<���m�|X[y/x7�Б��v!&��|g_�
�@��Qy�ys������.NX�<��oLÚ_ 2xZ��M�\h�����Ǐ�)��o�8n���tKD��-���x)!��B*i8�``9��[&`�m� f�w��|���+��η����,̪u�}�����ra��0�
N�F��rS�x㻏���ۧg�b���kfg�tվ���o^k̥��t�E���bx6�Y�չXn�����v��q�؅f��80�0�lZ�k��~�Xk����{�19�2��������bF� Z���8�x��#�������|��ް��?;7��.�!��%��-Oc��<ܱ�iV�:��b�VF�Έ'B��{��i��w�s6Rk��Jo�gA������w�wg�C����c����z�.����^��k�L�?������ۉ�X����c.ez��n^��F}@j�V
����Y,>���7�?c�H�����Ѡ�?O�Y�:�ef���k^<�*�-�3w��0n�,��VSo��>h����-�6fJq��6ߴך�%Q�d��6��eE���FIb�U�J�b�#也0?��sy���5�]E[��f��+�6@n,��pͪ>�wG���f�"�A3�����6A��n���킀�î���h���I]�5r�EN��H}��
���#�@�H~��Ԃ��	E>(�i�g� �ř=�th +��Bm-�D0ĮR�Z���dfy-X�b�} ��Y������(�������6��3�	`e���� 3�U&�a��+^⤿�ZY�,F�(w����(A{�)�3kL>��rxs�毠�:�����s7O'@��|!���~E޾|UVۃ��������@��1_��[9e���ǱXj�:V��N÷<����r�����<�;��H��M~�%���Ó��q[Y�����T��vm��p6���F��ƢҘi�{~�hCČ=. �O��:<�A�\�V֢n�7��Ѻh���k_� e�Z�\KE��C�[��x�A?A[�	j�`��!&��=���3�]��g��D+���B8d�t�.N��Ǹ&��ݜ�!�,`����I6@̧�Hd	�����5��9�#�Y��$*gv{�'F��OU���-
�@�\r!�Gq�U�`�X�r��k��7��.V��W@~�^~4�n�P�$�P�f�с��z8[�9��荿�S#�BDkgx��{���t�%{�W�r|�g�#'�[)��� c�����V�,��fB�P)G�� uk{��=O�B�l_�!־�9�|z��y����3�͟+F�?� ����I��)�H��[+�����u�T�-^���l��d�rGb�����h��.�Y��E��-�h%��?����������Xa����.ܢ �ug�A��ϝ�p
ww�I��F�о��j�%ZJ1����I8��܍p�eI1�Z��#S�����U�d�Y��n}E��;4�H� ��N�c�x���ZN���}�(��q�U��f%b8�YH˨�u�J���m�[-�)���2#�Ѐ��ߒf�H����%��Η�L�5-��[��%�3a�5Z���v�������}eG_*���
���ឞ�9��uo�csY��.����r���Ā-��)����TC�'af�9��¼
)t�����z]��疃-�3�T���jO%��g5�[+�7Q�BnÏ"�(�jm��mFu�D����/�P�k��o��am1�4K5?�����<G����>�`�o�;�{����#q�C8+W�����G�W���g�wJ�KgP��!�EK+L�Hw���U��y$%�?��ǀF�v�2��~���_Y�L��xX���4[�D�VD)���d�@�ޡ�:�' �s8���#�� ��>yE�lL�C7���n�!1A��iqM� f�'�A��]p�@�r��/->��
8�Rc��Qu�%�����ʀ�� ����*����(��o(�KX����f�׍r��nٜ�\�v��t��^j�/B�����N'e��@Zd�2�]��|�n7*<�}�����~��ڨ³TX��ͪs��'c_|Dfx9z��mhyl�q�4߾����Dlο�x2�_;�3�:�aZ�h5_N��e!����c�n�,�c���׿~�Rh�r�7�F�B�=�z�D�_��Y�
����j��-�f��j��^ˎ9o�Ǟ,^^�{���QFT1g�J���aG%h&���`�{��T�ޑ���J�ݭX��%Qvǳ���G�X���D��?��[��xj�g��� rGHy?9��d�59>}��ջ͛\{igL�>�����o2u��{��{��D�ͫ+�'�$����`Na���3~�m�=_�:��"˙xJ�6z�-��c��c��E��T2����b�cb$+������)�K�p������K�����t���{�K��6�j<odҺ�pcL7�d:�*�$��[��� \%�۩H��,���i�l�3]|�u؜�E�&_{o��=7�/k�.,�FN�J&¹w���T��S�7���.��[�ֱ��� ��H��˄t�-~���^���R|� J[2�)���sD����l*�0��{�r�	�Ok���͂�x�N�y�kڥ ���.��n}�`����8擪%d��ҳ��#�n֬���:��KY�k�m�J��|�)ИV���p�W'|r6j�ܰ��-��@�������_�y�k�Q}n��D�e��Qs�Y�Bwq��ʄ����a�Q��1��e�%^�7��X�.\�,��+
���{sHDa{Mn-�弋u�R�tK?S�	����������.e��v~��y��&���#P�Sv�E���2�=~U�l�W ^G��s��s�st�����q�{��Pc��n�҂Z������n���5#�S
��R�l��kƬ�Hr�\��dH[Ӗx�$\h��0��Ub�W c�ۺV��M�^K��*�!����U��)_�O̐�� ���c��1��'��ߩc�]K6l]�߮n����ӄl��YR�P����&B��\���m-o����Ѥ۩��, `m���QA��Y3G�gi=��N�	��ax��}�*Ϡ)�d��us�lT�}T��0�𧇝���yF����&��4�J����I>q�s����
�|)*�_��1��L��
5C����S++��A@�^M6ߍ'���u= <|}?l�?��2���kA��@@��A��	��������#�%��!�7���{��y�̞��^뎉k��%+�˔��~O�)���ǝ��6�l<t0r�+�߷�1������!����x؅|f֒�E
���~k��D9���s���^��v��	+
T*�M߁�OK*	F²|��E�l�@4�vq�σѷ�/�7N�S��xr�c����
�ڱ�����y1��`@�ڠ�L#�� ҃γo�7C��b�/#�{��Z
eE�XP�I�'�����{"�!O���3����'���f�+����u�AG�%^ڟ(����p1W������I�5/S�y=��Rl+���=�O���l�	�Yw���NR_7H��{с��f���NU����V�>�P�9��M����n���.}S#0������Fԏ���O��s
c�+�����r���l�]�L�~O,	���&�x��*H� c��,��3�G�bZ����g8^5+Ϙ���E��#lȽv_�T����^��~�����+�-0���Q�7�ߞ�xO#ş�*�KC��ߵQ��S	�������n�����s��k�WC����n�Qu����'��<��<��8q%<����8���=2㢎�6͔{D���������{O���j�N~8+&A<-��THC(��1I�,ޗ��6���\�KY-D���*V+�ϔ��)w��&*�dcC��.	;1ɐ���7�Hw�Կ�"�����y���|���Y����w'#�������˰9Q
e�xc��#��܈��@	A)%S�'����
�/������YY�͡��`���(,L�QR��?}����2��>(���h�Z��دE��f�Y:��=`�1����z`��o���������~bL����U���D�f��̇���og�~ʣ�5e����IjϤ'E�,#��8Q[D��G�g�%��|�E�P���A�^�mD�,{]��`�l)�*��5ě��e~:���xp�`@/0��}"�X���p�� ��.c�o��ַPi�݄尀Q�+pEQ��4DS��헊@<AF�{z�˲�����S� �;�I��\�5�:�~��b��@RK�5��"�!f�Bw��E���'��֏[�5�z�� ��*�`���гۅ��8���b���|����dI2��j3�:�����UW�7VQ�h8Da���d!��z�bJ6o�i��!�UzR���� [�R�,�TR�&7�'�1��N�������д��K���/�C�.˲�t!��������O)�py~�b��P��$�D)�@lgL��t������1�\����lf%��v�^�vNcJ����:�3XQ�8f7�oR �E� ��CZe�]/���Ջn}�uVxq{;+�GT��ơ��\ �����'S��k(r�T�� kt�o���^z��H9���}M��KB���󢾋|���o|�Kф�nWL���I�we$�?�E=L�;�E0��u�g?\R�B�MK)&C>v|;x�pf{JV3a��#
d�$$�(�;ﵡ��1�m���_C�|B��@D���(q��m���C�<�i��ls ?��1"���ps��zx�-�L�F��_?9��^�2�B��̭�ě���Yc������DԒ�/���t��ZU̶��<���W�����LE�@�ɯ.Gx�w�FZ5sW��|a���0~d��qd;:B>l���]�}}g���߆lϧ�s2�ԟ���Ņ�K�����X��an��^�P�9�s�1�De(���Բg�։���Q��Ӓ|�����%\�6�0Cάg�����B[QTI	�k䈰E߸ƾ��$>X͝W'����F��	j3���-	�u)~��Tr�	�I]��W��+�2���$E����2I��#��y?E��=�$,��
������{I��E� �*'�(|yxו�?����U#�Ub�H[g2��֠�uҏ!Jҋ����ˊMu��C�si����^�6���M�aB��_�+��|Ų;1W�g�D8;�0	�\m�5˪�[!i�2��1Q��z3��ׂ5�<�'�����T��58�+~�G�#�a�b�p1�;��������ڔ�����BX=��y6L��΍��o�!����b�J�g��艻�lL�����[�~ր��U�w��C{����U��b�T��g��1�Q���?qwrl׊�w�N���ץ*�%�b*��
��W"�z��	_��$w��6r��8��`�
��dմ"�y��sL���p��\�?b? ��esv��M��h�?eh_��C/4�hg2����M�ʻ�$�kG����.�I�{��l�=�Y��)�;�l|p���X�c���M�C򬂋b[��iĉ�D��s�l9��	k(l՘�X�,B;jӤ`|}�#���F9�`��D{G*�.p񲊶��
�jE@`�����F��Y8�1oL�b^%s>n��0.<`����+��*Ts� ��0%r`�MBJ��QR��1�����PZ��n&G\��+�-�3�����>�@�3qP������ٸ|��ע?�e�m3��Ԉ�b�*��I�����gu�&2�5�*�I�	{wp�����j'L棄d@<�����o��t[$�x���!�ˆ�E�9�Hy
@����j��=��]�-���e�gO�m�&k�7N�r$J�B���������:��;�[v�6��	>kn���u:"���=[�����d(Vܚx_�5j
�%��zr"�,���40��m���$�ɪ�@�����wA���K�\j�ʱZ.��i���iZ�2�ߕ�QbP`an�S=� ���=`�p�p�;��F�c<�5�(���	��1#7R��	���D`<�V��ٝ��-��S�%1�><# �lk`Q~S���⧰<�x��Ӊ��}8�*��6q//�Ð�D*Ck���uL�;�F���IJqh[cC�Ӽ�zB�b鳟�
���< ����(�	�'�Do�C�8�TqIc��Ʀ�U�$�����yC<?g����A𴆫��F��3a��  ���m�)�Q%g=E���~�jjq0� �6������i���h��^
+�fB�4OUqK��Q�5:��4�6f�7�>d�~�Kzߠ�SAK:��|B��>%�G� � G�`�t�� o����p?� ��Gtㆆ����:���{�Dַ�?#��d1^��HW[)�ť�F�<J���6���u�����RS���\�z
0k�珚Z@�zk1��"�h㥃�˸�y��%� 7sQ���;��Hgv	1x�5��ΞjԵbB�O��Ta3�.���I�3��z���)d|<v;j�g�}�.�fU�4�7P�`ӛ�[���P��s�;/�&�Vd÷�P����J�8��6�?Cb޽��=���>�
����%��{�����DUC.SZ& ��N�i�S፽�}z�qx[V��1�,�s�%^1��Д�����˭�Ow�'F��1�!;�hTվ�_�cKθ�*�;��j-��1��XB]#�E]O�t!;�좭��[/��j�M���x:��%j7[�%������T�V�p/�Z�#�ͫ`��(���Lc.�L�ڽ����a���ヸ�IT�,,�w����!����PK���#H?w���w.^��(v�&b�v���l����8�Hyذ^f���)5�gDf�%)???5��X���Or|����&�77���!�VڃQs���I�=d��]������]5Y��{Z� �����H��l/;n;�IN���]]#�J+�ZN��O<$�l���G�,��0+��4�m�p*��h��ѫm�0@rIlXx-�Dd��!�w�cӈ�O���t�'�����e�6c�9�Cf��3����*� ���p�W�P��׬�bN�[�)F�?���C@8}$�8�9����\b%H��=i��l�c�?Y~�p�|�i6��*���<h/��8�(����>�6�C�bF=Je/��~G/"`lח��:�%�f4@5�`�"f�������c�0K�>,�c��wM�W�� )@���Z���/I��X���7������'7b�x1m�D�H%�~n��4��vS�Lu�Z-��r��Ap&`��a��v��$6ǩ�kq���r��c��I�揸HT�ɉ�LC,���;�B�0O�����C@hi�fง�����0@~Nua����}�����E
�����@J;g�O_I���~���g֞�˰M�T��r&e+����i��z���|��܊p�~�`��ua& � ��G�u�SRh�Yq�
'��������p�>�Qx��M���]��^��P�rޫ�����+|xU�"$A �&�ْa�d��ݾ��-��|�)&�e�ܗ^�L=?C"�SB��v?cz�`} ����1�m{�#A�y��_��c��`�!)�MT)�y��W/ۗ�c���ԅ~��A�N�P��I�����	��Q�%(��Q	+d`?�決b��yWx �E�,&K��9x!�%l�ki����.���ڛ8����g��pԫۨ-yWg̵���'��6�_��b��L��ؑ6��a�P<$��F_��O/0\mP�B�����	к&�����Ap�}ɮ{���nʸ!�YTʝ�N��S���s���n��s�P�h'}4��nz���HR�}���;��A\��=!�Q3k�ڶɛЍ[���G���?�$]��#�Y���B�.��UN�����t\�U2,�Sd��.X	�����Px/Dz��� 2z����Y����w!����d�E���/ّ;\��6�(<w�+Ƣ�P)����c��Ó�F<���c�	2���jwfi�
���Xq�,q�I� ��®�fx�aa���d�yUoخ�Z�2�61؀�'���V��K V���պ��Y�$�c��AIX�k<�~@�����"5:ɑ`EP�H��t��7th+�)l�la�w �"�c� )��*�ByJ"M#�'2���bI����a ua���ꂋ(����#�0"�D�N�A������q�%���c	�p�_�ǅQ���"���HB�F��@�р�o�ʩC{�{�^�����OF��_K#��[��" �{�*�
�1�j<T�ԏ�39���'>8s4i}��n�hB�҇���#��o��ԣ3B:W�=#IG@C�j��0iX�'da��/?d��p�'��D���F�)Dt��ڧQQ��҅��	��~v�EcK`��zz��e$b�ěo�3'F&��t�	/���TH�8��Z&%�'�G��G�a�w�����+G�+k�Q�Ɠnh�"N�rR*�s���zh��	#ª<Ѽ���I.�QadY{l}�m�z|���~����>�������M��dj2��x8q��y�4O�(/�^ONJ-D�{�K�u�~�G:�obM�� F�5#nU3����X�U�?E���ntc�t���M�{�v2�����_j�D�iq������ݳ�{(��B���i+L�_�Wg�_�=���	��[g��]mCE�E�c����q�t���I?�J�Q:���Ј�ڋQG}��-�Ȳ}��(D+~��� ��2��n^px��:��}&\9���]�)R��g�iͥ�1k�,������G!�|��C�)�go���>\�}f�p4�U.L0f��'���`�Z6��$\�s	���I�?�o���pyr�W��.�|���}չu�`���4y����<�3���\��܊*�2���⧙����?П��1��?Z��uަC(����<��rr�SP^!h�����^��z����Go	��������xԟ�;��+`���qd$�W����v�0OPB�w�(#)J��:�O�����ZPQ]�>�r֩�v�'!<�����U+��r6��gg˾����;'NbR�iqrO
��I����ט�c��GV���v�o L��rT	�4�Ƌ��/��+���HK[kM����<�Ak]�?��_@��ŭ��1�xీ��XXX�<���E}�R����JQ~���P,Z1�B?�|!W�؞6��α��Ib��H�<(�������B�IS���T �K�_|_��ȑB񽱒;@租�"��r7�)���Cx�$����x�����+g�	��+e�@���"���jGפA紙�;]4]��!�����(M�zU�A�4����5[�☎rr-���Z8%+[�W%�S7ʋ;��/�lT�+]��;(zy���A�����j^AZ�j�� ���=rG��SB���Xcg�b~4�JZ�dԗ�<�$�r�8�d{�l:[�P�b�p
M,���!���ʕnR]��8Rb��h9~�4����r��N=�]�t�JU�)؏�fr������Սl����!E�"��B;q&�������Of	��F7AϏ#����'��)A0�
ȬD_��#� �J�p���,0�A�?da�4a��e����[��'�-���� �I�W\���ȁE���m���P�����9u�����Ӑ5:�P�`��2�R:��P[ �*���,����)9�$K�/{&��@�s5 A�U҅��!2���<�bl��g�3�3�чb@�t3æR�G���]�8���c��� �"�|���d���j�n�i�
+?�t�ń�tr�C�E�b	�(��Ki�*��6���pO�N�x��P�ި��u��:����󫌍)�m=�ġp�?��%35��l�������9��gw��g�ֹh(��	�����ų!��F�r6y��'��U:QqT#N3��g�r<��qY�'��J��#r��l���d$����e�c/:�E$r�"�'ԝ���_�J0�;��Qܸ�_�b���0���#d�_��J�kξ��AL��z�����/���N?��1Cv��3Z���{�"伱�w��K���B ���� Ka�Q��QG$2��v��}Dd=�/��a�@�����p�xK!��],/��*z��R�����'{���c03R8��Ԩ��}�	Ӣx��2�f���L`�?B}(�1�Gf0�ӊ��!���ЖN�B��d	"j	�!r��U;�B ��N-���֑1�"C]cƒo;�=�����Nt���d����)����Dli�q�]��]��q+�κ��d�~�b,70G=�/�ӊ:K�K���їc�U�Ց���%<^v
�F��kF����LY�
ǎY���Q��r��5_2��i�YB F����� ۓ�:p`N�
P7~�I�F�� �D����w���s����P��D���%3ih��a��8�n���!�cf��[�J�IK	S�gwke*���>6�m��ì���ik8�_pziy�"���N+ܯ�Ni'%By�����+?2z�Y���Ye�"J[L7U}2��Y�\,��Ɜ��z�P4,��qg.�̌I<����b�#��G<��rn����,*2?������g�|�����h�i�k�pf�D4����]ǭ�P_�<C��
���9�o��T��3 ׵8F(��^|�b�<�C*--6�\�C0fQ�[���N��@3�'Vn�E��8e�x�a]~-��+[_*�}O}�.m�B��]��Z�o6�E��Y�R�:�h�a�ah�rч�㯕׏S^���4��#��#+:˲bE⍋��Z1��~�Fd#r�C�� J��5����R�P(�=~��x����"
G�~G��!c��2���f�?��:�p�OT�1T��8��9�S(Ҥ8�ڊ�I�E�N'�0PA���%E���nE8Fsap�ԅ����i���-�ɛ]��?& �H���1x��U؀�@:d@C	��a�]U܉S���Rވ�xƣ�������VYh��3,AV�,�� I��D���BE�6M\94����a�4X׼���M��ו�����	܇�Y[tO}|��ss5���`lo�M�PsEg�����6�[�9��i_����s E'�7���ui���=R�����ͧI#��ށ��G��P!/K�zq� �a��[Fa��4�%����C��b�3K�@��0��	k����a�ۯ�4�D�Ί�\>���ܟ�z��	P]�
N��=LhS5����ӄ�*�����8
�cgb�XC��R��t�����s�:f}MU�4l�$Ż�v�;NG�@�g��`։�N=�z/�[��|����G�Wk��DT$��E"Hrthy��h�P�~�<g�����a����js@˿���������Y����o��f�];�v,پB���7b� ��O2"ywRD��T}2,���_����,J�=G��m=Y�.�@z'$&��1�i���>Ӫ��"E��ປ�"_�#�����˥��N%:M�c�����W!�R%�����v?��Y\(n�L�p���X���Pl[m~�S�~R�pڞ&�D�rG�Ul�O�F(w�3�<Ί��q���F��4v�xp|�$EŘ|b�ð�P��V"�5MC�PiIxY�+�j���;r� �oEY��9�����
f��v!�i�?�]�s�PH�P�by�Ά�:'���H�vn|�x�����u�ړ=^9��*ئ��E|���:��(��N��V2��Bmȼ�,�=��g����s��y\Q��dB�@��lXG�'B��54��eN���IT)��T���GW폏L7�M�t9�!�?��0P���B5P�n������v�]��B䩊�u,��O�Q|�Y>h%D�e�=?��CI[,v4��+���1f�(���� L�*��3 ��n�P��}�-nJ�T��\g�����s.Pq��il'�|{П����P\�qwU��Q,�4�&��+Y�^0C��O�6c��mՍ�ӭ����t=[-�1�b(�jD�t�';�_@�g��z�wgA
���S��+��1�p��Z��_�@����b�X[�ZF���(d��A&�y��;���Ϫ��aB���J�z,T"���z/[7Xf�����$ʹ#�s�O�'�<�����Dobœ���,�Gq[1E����М��}�Y���b�w��h�����3g�9g9�W���P2��E+�̝ ��X�"6]�(�ce{�S�*���P�`���f��6�e�y��b���>�!i���<������Kǂ%�nk����k��%ڿ̄Xkl�|�uMrQ���O����S��A��l�AMA�p��vi'w�B�����n���ڢt��+� ��|�0�u@Y���@�ښb1���P~��|}4��H��({����Q�	�V�t��
fnv�k��LW]N����@zU�A<������M�j���k1�� �`�Zʴv0ԟ��#�<\�c��Gw[QO��T|����D��W��S�Rڅ�ޔ9�4CJ6R��p�2��>✝����S��lG^�	;�z۴ �}%�V���_�c<8�`@1��K����c���p[��K3��W%mX���T�_q�H�Q��j��'Q,���Z8D���:�V~%���s|5F-g�mL�n�ɎR\`q�, :o7*�1�V	�M�"C�����������cqq�u�l�"NBP&ʒ�#hM,�آ*���n�`�g���D�3���?Ύ �=�}��ɕ�&	 ��5��f���vH�X:M)�P��kcV@}�e6"F���#�A�J��3\p����f�K�=7�m�h
����Z�T��ΔC���݅B*׋'�D�	O7 �S�I�K�w��3�w�މ��2/��*nj<�,'2�mr>���.�	BC��Ѫ*�\��2C�ƈ�9��G{Cj�2 �ֺꚄ_�W�R&7aS[���#�'ԧ�9�V�F���bc�e;�������bb��ss�2ވZ�e���|���Y}̛ܣ��)S#�OX��Kf*�B����H����E��6[q���v�w�|��*�ޮ��v��>�2]�*��4^f�S��w�a�;����u�+�Y�����*�43��&t@K��7�#���[���U��ԭ5�P�	��j�H�k���Um�\�%ߟ���p�6��1�7�7�Eo�Z��b�i�@���o]z�?��v����>��m���ֺ3�D+$��K�7	��U!M'�НPYBvyS�T�{4��#S'���YA[wcK�lN��$iJ<iѳ�(,	*q�	�	q�K�P;�	��Gő�a���Dh�N(E8��;��5,l!�䜬E�I�Ƌ,wal�ȒL!��O�hZ��9���h�_��%b߻�����P��N/tF�QE���Q����Pv�q��Ec�S��^�uI&��Ӎ��C��B��R4-&������|H��eDf�bX*�|i��{fS�~y���fT�a�*��h����9G�8�^�����4��F���t�,�����4��t�#���qzx��l�@�@G�̍�Q\��!9�
��r/WW	���thv쎚.������?D��B� ����nI-�NS5g�-��P�8�73D����[���7R�.��T7o�(s�� ����%P�y��eQ����.�!1@�>d��x#Y���沁 m�/-	9�_�Z�j�+��B\YDw�ی��1W��F/a��v�&ˊQ)ׂ1G���[\
H��w��]휨}�o�,jO��'&)F�X�K�y�TȁC��B��7μ6�� G�J��H18F,i$z�~��':��U�%�Y>��-7�v�O�!�� �ko�ftwa��"�p��Y�Ň���;d|l�zX��-Ck����|җ���F�5�7�+�;��	GMT�m��je!+#\@��e3D{c�����2Z
ϵB�����ܵ�c�{[>��9�4� �P�p�`��>����ԊЅr`4g{����x&�ez�jǎ�pΗ1�4�G��΂}�F[� G��o���$wC�Ǵ7��C�.�:
��=͙+��*��!�� �<�X�,M<��:��s���h����m���GF�<�]e8)����Vh}�y�a�W3Y	'2����"u$B
��I�p͏�j�حГ�9"R���*�s�o�t���	���Q[����r~�җF��,|�O.����S����#�nt�,�I��
L\D��mE�@s��.�����>��[K}r~1���y�����a7΍e85�"���!��Z��\�s��C?�&�g��5JQɎ����^7�1H���4Fj�y������c�Hq��d�Ta���[�Z�|�1�v�������fnl�ݠ�7>V���%������Za�}jl�ME�����P��*�u��t���(��w��u�4�㸱�mJ"�bÛF!w�7\��
兔��y��X��P��Uv)/�]�%;p`Mǉ�Y���X67��0�hY�W��%��<��~A��2�)�X�l20�刋3Ut�<(H��Ҡ���$�"�Np5��w����p�9eq�ɜ����"M�5Mo�Ԩ�Q�I4�RO��;A� ��=%�Run�+���[���RP��t�Z�W{��I�JՑ�1N�P�H��� ��ի��g�Pԡ�i�k¿V�.z�h=�ٍ�چO��Is�3;S��Tn�i��{'��3!�(�Պ'3�K��)R3;gC����'e+�,����v/[}ɞ��nDvic�m1u�ijV1���sڟ͝o���3T-�8��O�2 t��h޿�B�1�8� 쪙(1rт�z�!f�+Fߨ�+[1'�T��D夰K���R1u��*�H�I���.�C�7{rf���
���S��nӵQYX7K��*8E��N��c�B����͸o-?L��R�ju�R��Y�=(�w¨.���g��Dg��}�}�D�,��^��c�����#�q[J��t� )g���[Ȓ��!�c�L���:�O��:Y���PO/�f����Le��Gڬom6y}��Kk60�i[L�VЩo�9�UҒNp�-�I�v�dyj[>��VR�Ww0I���.�{�R����l؍U�2xrd5���kRZ���g��$0eKv����
��m���mO`���qT�;(������<dت�!LY���%Fr��&���R
�4 �U'���NHT�v�#G �s��U�%r�����U��4;\)�i��,��%�SU�A�^C�ƹ�F�Ҡ����J%n:��T�d!1v����[Ǎ��B���nU��7��ˋ�84�" ��o�/���כ����a���I�T�������]��	&��w4�V]r�E?� q-��9A��(%**/����C{9��Eg�ߝ�n:������sbAIt6X}ņ�O��]�P�*b�~�Ä~!J���<_�u�{�V��:�7��w:�7�<�S�le`�c�@R�vv�I'�ڵ�O���jgn���`�W�<��	y��eV<H���W�]���mW,�W�� �y8c��`ǰ/�=������۵��,M��4�Sߟ�42_�U�v����V޳�W�0���M�1��Vg�ȳ+��3���oݴ���?r2���A`�������d��C�U�)�����J*��N�]`�a�P�'K}�W�q��J��/i�Æ!��s���<3��`-fq�	ݺ�u]u�R�b6
�o��f	]��a����R%�7�.9����}��s}p�Z��7�W:����s��*f�O\σ���<2�\�_K�|L�I����ʫ������,�͆1�|2����ѼTKx{�ev�Ac��>o��q!	e�_�TN�K"�T/�!��4����:��8,�]^����:�*�V����jm�r�/�Lxض��/�D�0���8���ٺ×9e7��5�m�
+��,:��(�U����K���t¸٘�î��l+���]��ݼ2�j��19�2�65��g�-be>Z}�k�����)�}g�<`�)�Tm��|�{5Es���17�k����D��ωh�_-�l*.�N�Q'q�נ��x1��7�ۇ�C��G�y*�V��a�ڞ��li�_�X�	�����/�66T�I��It�����>�y]'S���Ph���}'ZJ������@�Sn,��%�0xt�C����=A<��f���v:���$���"c����m�ۡ��.2Y	���5�N5�_�K!Z:r�������������Ck_7}�V,q�o�)���):��O?3;��
hd�eXf��"N-/�:��9G�z[�����\��/��Ԗ�x)�{�ޏ`�
ɝ`�R�D
�W����`��w�E���&����_U��JG��h���t�卯y�������h&ݤ����J�_XlB�nr)z/&KSqF�~0/�}��m,�+��AU���^[{+��ȼ�26l��pOe�V�/�;(N���ɠ�+��Cf�*|ܯ��w�-��,	����@^��00�l��4,�p���z�DN�ۻ;��μΣ����C$8`���Ytl�{(M�.��+>���Ma*��1јy3�=�얍Q8�\&n�w5�@�V�lf������VH+��nq;��2��2B
ͥ{������_X]��=Nl�,���>�1V�qb�)y�u���V2�&��3z+����#F)�B�(�W�y�f�EKK�|x�Vp¥��4|B�Q���!O�:��7��U>&��F�z�G�F�%�+���[�#8����w��}f$��j㛑�ؼ�D�ovP�ٶ��j�>7����ƦD�YFQ���Y=p݌c����m�$)�B(�����h��*�ޱ���	@=�K ���۠鱛T\,z�	���lc<��ً��iZ�7A��:�g~Ǭ�NZ�?�2u��������=��t�O3/��hd�_	�~a���_d�2��!��V�ۧ��m�|�d�i����1 �:;'���\؉�U�U��
�������^�U�y%�QmR�ϫ��T�|9�Zޠ�U���e0J��4�k�k|�����l��7Q+��N'V�nvpG�h���ݩ�����
1�#�����9�r���Y��b�iutn%sV��ls��~�?�>��']�ZA��P�]��ƕ\���\��p��,�H����%��_�'�DKɵ���Pr9lto�����R���7��r�Xz����R���0Ҕ�e$���n	�̐
Xk{��u,�y;�Z�J�y���5�l�vB�&��_ݭ�^<�����L�����V^J��JV�e��#�<�
M=�;h���6�q�)�z8���k�;P��'����+���ZV9���)�ĈT�Mö�9�)q�=J՞Q�j�̠>7�_�צ]^�^��W�_�����d��q8^�����iu�>e�y�b0Y�t۷�Kd��z�rϿ�U���7��7����!�s���`nw�j��m��^l
t�딼Ѩ�v�
	n5�<>;��eD�O�M�_?�}�PQ���$O�ۦ��.V]���9����cd�^~�����gsԛ=}��#a�&��Y��~o�5n�oj����S�T���:��q$��d?�7R`�VW�1y9g䵠\�"�����kO|޶�Ds/�D���ǘ�>��G�E�{Q���o)�:4�PM--���w��][:�\ɉ��AJcJ���at�`m���Z@�'����9�����4t��a��R��1UwU�X邽rU|����&�����_�˫5BLKo5&��v��P�K�̋���N��I�MJX���]���"��<�<%�?T$���;ۻ���@țB�TR����k�}1���d��Q5�$ܲ|������h��cm�*ɳ��c����{�.POgʏ�+�e�{��Q�|��n5��,J���6��}��#k�飴ĥ���<*ܬXd#�Kx���
ڱ���pę��奸�^��.�'z>6�/��ؤ�誫I���jd��9\q�So�5�/�%5��&�Q�
1���7WkI��j�?[f���0��}w�˰ ���}9sz�_��p��m�}�;f��FN8ҧ6��������1����Cԁ���o.B�kzy�1�����A���N
��s�?�k2�����=->k}XZ"FL/�8Z"�}Q-� N^��~R����w?T�)����6��&v��ر[���n
�/*=|�Pv��U�r���dvi}ֺt�/S|_�P;*l�M�~�K���)zSnQ��̅�T���J'km�޻� �����}�k�p*���,�G��Ǡf\������q�m���/��%�h}�i"�^�-wK-�$�7����8��hx}��xxTS��\�����5��&�u�_
1S������%~��'(_��$Q��j�J{�S9���a6�E��jr����BX��>�����m����Y(�y۾ۿ����q�*�vv=��Lܾ�����.���	U��LIv$vQ�y��0�.��j1Y�ᨵl�!���p�H�Ԏ�i�ͫ<�����,�fnm=)�8�8�qj���<��T�W!��|%����3������{��b���K�әNo$���`[��	�ee��wQ�9{N�u��-��I��|���56|�>tL]O��A�8�K�L�ϖ��'�F��sQE�;�Αz7g�dI@�^���~_[�b
Nt����ں*הg�*?a��3BT.־!_h�m'0��W�Pxr3>�!8���B���.��(�t
G�~��kI�W� ߟm�|��gmK�P��xzѫ<ل�tU'�3�,e�ǉ5���i����oZ�sJe��,���\�׵a�ow�꓿،���P�E��Ng��9�����ԃq�\�߷ʨ=������o$��N^ر�#Y���5�=,�4;-V��<��f(_'��D}�4W�'�#e�{��^���c��������eמ���ɁY��i'.ċ�\:�޻���o��nͲ'r��<. 9����?�YD � A��1G��T�*,b����ۊs^ěSLW�����p��5��Lk���w_�ʋ3�/�=�8c��V=��nuz~�b������;��ّ\m�:G{:b���3x��D�5`q����MT��(rahr?��o$f�E�z���셷!��'��^ �T�s��g��~v=��
��θĬmu�M�YR��s7f\���s���,���[���s���q����(�J�)æiaR�l��q02�߅P�P�3�8Iq	�D���`0����դEsa�,�	Uwk>��G}q�)׽��~�.a���:��ݮb��bS7�Q��oxص��11P��:��5�w�k����ٺK��t��ZB��� ��ZP��@�姪ѽvl��Ht��-�!��Z�s`9R����lfrJ{0�j��+��9�P��8Ύ|�;�t��ɝ&��zR�,�^��6'p�/F�,a0j�y�)��y�h���`���t))ϼ���F�ըc��+x�v,�`��Ѧ��'���Ul�����'���nDY�,��#Z9�3��>{٥Wy_Iya�rz\�S�2���vE-���VO����U��~�9V���r��|�@����~����A���b?o6'M�~��J �O�J��̦7:����A2��'6C�q麍��C��u'ɵ�j��zG�n�� �6��V���z-�g{����m�_��.v�{����N�H7���B����I���<��q��o	<̰���m!B*v]5vFg�
�ݩ[�\v���il�1'�m��Ķm'L�dbsb۶�Ll۶�~��]�5�T�ڵO�9O��>A�O-Fꯟ�
��Pq�5�1O��s<��;O��O`5�hk�M�c��ۃ�I�P��y�&�^�������D-�;n$%7��f�B��)��"2n33��2ը��k����+?N]Hg�x��Նޥ���Y����������3B�'l�f��d$���-~��ȉ��d�y�\�٫褸��x���	��BX�]�J��6~x�Ѷ�g�pV�i��I���-u�E��C�^Z퍺cRIK:�o�u�"4�����Wr ǂl�).1$k���(��x�A���`���?��d�FF�Ǘ���,�<�;/ڦV�`��XB��a-��0���Z��Q�� a�8X��V0��
���MI-�t׸A����-^�e�D��߇|agm�^��Y�47��~�G�W�s��7U�t����'�	�!ϳq�`s��ZwJ+��,���N�C�A>B���"J��}^%�\/�� �P8�)D��P����M�r}�����:h	����QxY��ee^�0�ǅMfMU���i��C\��������L�D����y�(v���ġu;�� �RL�_���r�W���v�Ƅ�Xy�=���ǀy U�%Tv0����J�7uqт������q��T����ӦNx��~4֨	�:����{y��5�P;b��0�����ʄ���O��awϵ���nB����#6*��l��nӑ�&��çbG�fMEf��S�W�x4{p�Qs_�����1}�=�G@� ���6�z���q?ivKU��R��o�/�{'���@��u?�3;i'�/Sgύ�b��e�s����ٱiC�݀J�_f�S~�G��/��v�P'{��uM�BUD7�U�r������b����e?��	s�+� Ғ�t�Z���̀��^�����A>��)/ţ����.}��}!�ƹ��~T�HL�����әÅ;1� ��n�GR#0�tH�*Ii-��^��h�l6��}K��\�01׮���]^��}����C0c��7��0qS�qE|�t1�)��xn�����w�/������}LT󪯃��𢡐���:R2�,�\ۯ\���������t<��_��9���ӸD��yw��@��@�L�_��FC�v}�j�Ϳ�")�y
@{A�:����ҼO!��0��b�>70k�W�6�ɛ�V�3��)E���~�n��?�rf�~4�B��
vxmo�'����,����я0;HD�/����$J.Ns<��\p�'���E�� ��&�����Px9TtݨL�*�<o#��%G�a��nփo��{8�o��3�>D�� ލ�V[�f��>�N<������ImŐ0��焆�k*9<%W���H��y|O����؇�T~||�Ȕ��32m���{��/hkC���u�� 4�WۆT�t8T�G����%�	����R��IbJ�r�̌W�-o#����H��w_�1~��Ls��<��x�R�1$)m������@	�4:	۱���Ki��/˨���ьX�6�Q��.(�t��ic�k����3��)����ρ#"8��tC�]�6�j��6�xk,_r;�[�`�������������d��֣VP=1$Y��#�r81br��"y�jr��A�SEQ��?-?D�D���	�d���*h	��^��ơ��������<w����Ui+Y�63�}��y�e~>v$>���2n��.���L6���2T�G0j=�q�N@tא�IV�4����i-e��&f�{�K"j|�)��Nx_�ٻv�\/�Oa�S�4�,10� �#�*��P���I����j�P�xi`~�%*��J���98A�Ο�����jjw������#��vI�\��dNG �+���U�M	�H!����V��{.��4BH�E�W�`��nn{F6[�<:��r��]�w���5*�wۤ�Ùn�ō�x+p�R]�ݚ(z�นW{
�0�:�՞o�?�h���D���T΋F���k��#�כ�p�%�ո�0*:9O���t6~�f���d�(ȑ��;KU��G�3#�خH��5;9ib�X�5"2�[Ȍ��i�[>N��/�H��ę��m��|�!�[�7��0����|&y��vҢ�3� ���8�aj�rM�	�{�g'#���C4Q�EV`�G�.�����_	!��?�6.c0�ŧ�2s-�Q��bl�h�zs�T�!
;jK���x��s6�_���E���b�I���#��̘��=��z���I��1�ѿ7����sU�����e6@M���7j��P��'��G��o��2��,��f�lDZ����t,L��M��6&*{Kubkl>��)4�ƞZ+����{ ���s���-MY�ͯ߻^�\���C*�4�H������&j�b���KV���ņ���U����F1��<������u�o�� ɖ�y�W��K�
�N��ĤJ����UZ�S�IAG �Ҝ��Ŵ�*�5�n��~:X�C%�a���K� �+�?�/=KSá-&$;��,�B�ߓg&�f�	{�PpUxk)�o�e�8:��"I��Z`�$�n�M��@P��~�[�U+3y�ŴA��Y�+R0��CI�Y���Ce�t��?��
�{�Nd�mw[�ᙕ����b^zD�/%���'
e]�,� ��l�b��0W�I�PeQ?����a���$i&�G�zr�	�����p�x��㏱~Cّo���F�J����;�i2[Y_XV*O���T�+�C����J�
��rW�,�$O��8"��8&���a��˗�\�<\�F����n�t��W�1�����s\|i����EZ
4��d�PY�7.�Q$��%W��֟3W1��:P�o\Xl=\�ۣ���V��(�+���t��f� !�2�i��R3�|�X���U��'8�]�,\Yt��¤zEX�/E���=�-ti�)�?��G�gL��ᦪ�z����	&C9�Ȟ+��_�ہ���{�v	�諈�/e.�?(@�P>`8s�������:���5��^�w�Ϩ�woj��Ո�$��~g0��4FX�@�;����)�0L�Dz� UC�6G����̰�T^��p���`UAP��GL��e��d���y+��X#�شR����a'��ţ����Ԥ�B�R�S��3H��h���l�I��1n��1S@PGlG?t�{�r�����k�Sg���(G�=�sHf&��=�.��"ҫi���'O����� E �W6f�j�yĩ�J>L��a� +#�6���!��)�ݚr���U�p�%{dj�&�̍ͬ�B�#���u��,M�H\-<IHq�9!������%)��}�Iwb�.�g+:�Z�&3�2$ LT���-Ѩk��J'��w���\%)��}�r�����^Z��$�>��c��4G<0DZz�Z�R?�Ecil��o!��	�@�,��;�i<�2�TƏ`���3#(��0��y����OJR�_�G�MS����
+�bw����X�R�I=,��'o�Ȏ�3�ϟd���5�4l����1R�S�Ll>�?� 1�mu�32���N6�N�us3>�l�Q&�d��,�A��	3�V��a��a�^�iz�XL �,?�T��C�������<=!4�=TNX� �]A��n�@h�v��ڠz�3q�p��L�TN�@c�?�a���C���lH����$e�Ml�E���!�<�%e�Ϛ�>�M$D<�(M"	^;���<]A��8�K�����@0z��nx����$�b�g>�_����6$��]�A�"��fx������Mb���|��c�p���aVꡀ��Q�Q$�c��ʇ�%u#�,��?�
�Ëe�qS�������Zq����EĶ���~}c��6Q�l.Xp7H�^�܌�:�#7嘭���{��&�~��k~�:P��bц�SX=0�A)IߡJ�Y.!���EZo���N�K���cMoS�8���NE	f;&KF��.ֆ��O��(l���LUY}�Ø�}5�Q)�$�<����5d��xE꿯R�q��0��䘉W��?Z�z�j�v���c���dzl8��y>]�=�/�g�m�Me�Kfz��ޭ/N �d�3�$�s%�N>�Ǿ�3�(�%��(j���� ���3T�[)�+~��������HSқ/�#i�P(��L�t�Tk�*E®�A<��bsY��&Utq/���ѵ�f�Ϭ.�ׂڣQ�le9ڭ[d�+:�}�R2	��03��~�6������]xf�W �[����o���?�Q[�����ɔ��g? ͬ!��3�͙H��?FsT(��Qq�]�*�9�|ߏ;���?�+�����dc^�>�z��.�FC���r�"�g������6���d�O��zo
��w��x� U
�ޔ�1!�]3%���m��0ah̭��JiLշ�J4+���҈�! %'�٘��FyR���&��T1V67O����J�J��A� �W��Dhg�KCvy��i�
܎ 73+}����Ji�,A�e5`�Հ���`�{�]Q!����_5TT���3O�<����G����e?Vp�����v����?O�d�u*�b�"6�y���迚��bF�M~�i�cUA��:�H��H�e)ju�-���l�N��:����Se�)����	���2�|CQ����)9�h�:����T1��p���UR�0��R���+-g��qj�R��<l� �/��Y��:�k�#�
-���zep�����,�ཅ��Y�+��)��m����;:�9�N�Q�х,l��������<Bs�a���䳩[}c���0jq����Ԋ��$�l*
�qIy6�A�I�DpY�]��VMU�jH��y�����T˂�M��z�4�5	��(�+��/b���r���k�Yen`36��]�S�s�l���Z	��;M<b8�^�����:iKzK�������E��_
Gu�;�a���z����N
��b���R���"8�m" ���:Lk�/۠���Q:�d���8�@���p�<���� k�e#KW�,9��?�|)��.i�涆x�Ϻ���[V�	�|xY��u����Z��`]��	���L6�ͫ��1�"���I�e]
�`�a3�ݟ�j���|�ɿ�[=��̲s���Ŵ��X*6Q[��N�]oX�y
�=}'1	~�*������ᐪ��TCB�
l�4��C��U�n���/����$�P$i����s�\aĻ��@O�]�4�<���n�]g�����"�,��􎾸���%KHKzM���J�t��C_V��t(d�s���fC����N��$s����ك<C���p�1�Y�"9��t���G"�ٴ�{7�|���N󙾂F́e�~��)�R<@�ݡ��-��F�g�(T�R�EN:%[��hK�@۩�jQx0:��lMJ��i=p��}n~fu:��I�G�gtzK�&��2[��cݺ�$���m4m3���ڸ��|�����~���1b�$��?~bXmMQ�Ծޅ��Y�L�?����� AI6����˥Y�M�鏀ê�_�(jQ�,���q�.`�Z����2k7^�;8��g�jy�}w	Q���'g|��C���8��l��'X���P��C��}K��ץ���ʒ��Oq����Ҥ]"?�]���B���n��y�7�t�>;?d�r5�ѳ-x𝡣��5�:�s U��[|���<z7�	��՛�
*����]�����ew ���ѭ�Y6��?F��)u5�-S��^�ɞǿ)6����DD�nNdU������@d��_j$�m���r�����Қ4�f��J��ٙ���<�$�۱n%6��r\�9���oQ�����~k��V��5���H�)�\>��C%�P��:����Ή��#Y��L������Xw-	���Y���6��Ū�}���jf��a&�\4�_�΃��m�=�����S-�W�ƙ-�v���
>��q�퐖:�=�����JM�:�jx���뫗���"��Ø�B��1�3\&bh��{Q�Xr�gV.d���Tр[�Q��L��\~Y_s�����K-���t�fKD�jAI�����]o�?��_k�,r�ĝ��n�.CL�f�Mhj}hWf�m�N��-Y
�m�����j�g��;
��8rs
�_��ni#:`��?[�	�k�~�09��<����uO�'MV�~��N���HZ���ܷ�I<mc*O
�V��Y��dI4}b��2{�s��W������.<6�����Di��p���I����$���-����{
������:0�@��a�L�)p�bRd}���������`��KC%�p��.�7V�Q�����_�a�/O�wr�4hW޲t~�}��mD�!~�މ�T%Y$Z�G�K{��+�ӚN����N�d��L+rR�Bc�JP/
�G~�ѱnm|��w��
�]+����ߨ\�rn)�$�5��=��˯���T�B.+ߡ�p��� ��d�äF��e����:��94j׷�6�;���9s�z��=LA]�ͫo��Lμ��l~�K#��ށS��|�	��:wi�;M4.�#n�����������a�X�9SXd�=��!=4�r�ĸ����S`6���]�I6��}�U>?i�� �.o~��Y���_��0�-x���#�!��m�x����hVڸ]H�������ǁ�������^�j�lo�[7����;#I2/���%�J��%��Q����2L�qs�8�G�����G�账z )q=>��a��8�߿t��W�O�zh��"���M�E��N�ꐷƃx�vS2d�?O�&����:Y��>�(b���؞��`f{�<���ڄyJ���S��s��p�a�>�ǂۑ�>��;����87m]�d��9g�7�ӏ���y�ߘ��I��d�(f�n\x'''TRz��]�X�%té��h��0��y��)��������ۧoB{�c�Bq���w8��sTs'�Ș��]e�<�3_�=�+x��А��Ԗi��Yu9�ǈ?���¥dX±����;�����}�P;C��B0�8P��ĉ��gB�au���X(̴yƐ��Z?Wӛ��������r�,C*2,�$Xa/��v ��4�>},�F�]�u+>�������;�p9�l#�	FЀ���c�A�_�`�o"�
�S��oC�V�sb��`���h����Y�PĪԪ���Ӂ��.p)6(c��S�}�h�� �o�
l�W<�{��vkFN�0���4��R>�Ĕpt�_�w�;l&��$ VVd6���A�E礱�N͹:-��܇��^��:P�m�Ԣ����"Z�7W(?�'�=��*�Kۤ�dY)�V�sO���F#Q��.��=�%;����R�&i��ԙn�{���@C���N�-c��c�I�>Wq�E�-ة�����g����Z�{�VL$�����]~[�@Z�Q�v��t�L��d훠-X�0f�/��]�)s7�2]�QB	�m߱]�1�{��/����<�as�!��i���]�mN�nR�ṅsV�zk�̛d�X�1?@~�0\�?�=��&e��Q�o�,w1�7�no�e��
��{gH7�ІVwBj]�I2n���t>zA������_��"r�l��oc>�ܿ�0d��甩�Xzx����V����줛Wo��(������4wrv��E���6j�HHS�{a����~%Y�����Ue����Z��&U��l�;*�dw�~�3�.�j�2$]�~��nA���������}�l��0^.V�a%xEpY��t��Kp��t۞�b�w��"�`t]�(唉���ʔS�]�w��l���/(��L"'w!��#"�=��/a�*R��i���#:��HV]���ʗ����^�OM&��w{;�i|��h0d�!��>�{����d� i�Iuxqn[�W����'OQ7�jH�H|Tn��Bi���Ǡ�-g�E��q����ll�8z�E���2�
�Vc>3����pW^���5�"���� E�ݻ/��=McU�zM�VI&R�M6�F�u�C�g�mmd`�~B��^<`�����<i/*<��q.{J%�3t%�@�2�D���]X��־5��e��=+ι�w�/�!l�3�\���B�`>f��W��$3朮�{���J����n�z��F�	��l�h!aXw
YI�|Ζ<�)'�M���tEFP}J�܅I�{q�(���eV&*7u`n�����;}�8G$�E��
fIɏ���%\~" "r�v��נ��'8��I�I 55+�Ļهc�m�/���k,T�9:��� ��9�d��Yհ�i$���-N�5QӋ��B!�iz<)sR���� ��ߟC�%���ZyO���Ä:!�V�޴M�A���n�"��X�xdhF�r��P�[�9�0�
v�1R�a�qԀ�H���2��w^��~4�v�#-�Bڅ1�@#�&7FRa�]�๻�IxZ��w�G�ʾ��M,� XY�F��8ث�f�;�s�򥓴~	��o�-i߉�؏4݄B��`[�Ļ8źՀ&r7(��|[����A�5�6DV�U�l\� � ]�jj>��"r,a��z4��$��
ٿab�e,�W565��(���������2�3��ow�R!�j�KL���&A����KО��O�s�e���R��z�	������n��}�;;�E�cn��ꊷ�\--jڿn3x�WR4��:k	��B�9Y`���S׏�o�G�ѥ��Ħ��V-������w����b3?2+0�z��
��c;$�.e�"P#?r���B	,��X5?�����]�y'�NG�XŎ�eɇ��y����Vۿ@��9��NOC2K./[��(�O�b��4\� ��tFX��uq��G�H�n,�8x�H,�ϙ=�O���EIv����%C�
0y�����N&Fd�Vk�����֗����S>>_'��B~�[_��TM��CW1xZ�D2I�B��Ȗ����0QTj^�;�)Ǳw#���Ŧ]�]��S+٨nuTL�7�X�qO�eF��!���7��y��ײz~�8-�N��g&z\���_>�c�	���	����!����њ�X��-+��l�S��I�R��5�D��!�ȺQ�B^�s���i��g<Ef��=���T�d��|4cw�`A�%�ϣF�bHA���݅n@�uD>��=��J�7eiǕF�7A4�+���xu�W���a��[e�7X���3�+c�'E�X��@_(��.%���s=3i7�A
JLh2�}�����q{�C���̷Ov�Kr�q�)��գ�	uX���y�NRF-ր�_:H�B�J���ɯ�����rj�L���y�d-'T�C'W�(>t�$��� �ȌR�hs�T��/�)�����%��Չ�{���fq7l��g(p��o�Cb!#y642hwY�2J8�6���.R����������V�S�o�/��S��� >,6�bra���"���i $j��BJ������������e�a�x�-��0��3攐�a �;^F��C	��Y�Lg�U��ӵ4|�>-xM2}�J�01.3�sy#����n�~e������CFS!���e�F���i;-��]�賫=n�01ɚ{HL߅�� �UT�쁶V�ܢ\�m�y)h|)9��k)����ߗbo�f��E��5��n��L�Z�
!fɃ�=�9�@������Ҏ����m��+��<���b�r_��r�M#S� ��h�����
��{0*bM��P��C&���<oΠ����g��Ub�8���C
�i�(ad)��
����$�V�$�NM<��$_���0���.F}6��W���@BX�k�E���e��u1��"SĞAh"9봢4�/��~r�+}�����e�`o/��q����M؏9���ȑ�?��0i]� �nS����K=����Yt:�Q�n���OPܓ�lX�gٱ��z�aAP���`�fݴ��ZE��aȸ��Z�4��N�xsp����*��a������!�i1�v�C�'8�cI�ѹi;a���V��n�.�f�5�q�Agd,��(c�:Ȥ���-��O=Se�D��>^��F���C����w{������~�fb*R/�f4���\�71�J�3[��m���ܙ���`��,��U�O����
��7|�Bp�����?v/�9ő�������*��~�� ��N6�IT�3�h�(5�Fvd�m�	wO<�*&Q^zמ��!��������E�(0���D�O��I_�Ļ�7/vH�!�;�����ń�������`��� �7��qхˇ���]���LGĄ"R�mT��f��}����n���z���h�ah0q��+4����^v���s-Qُe��ꀦU�j���&�[ԁUP��g���I;.�Q�K;pL�����w��3�f��A�$��z�m�[�����Ш���C|�����6G��Qq�䧆 �Z�~!P�J.Mg�zӅ#��^��;�H-�u��V�V;���{e�%Βa�"��������*kh�s8�V��U��FV����z��N2��ee���ݲ�-B0� ��&�uv�F�D"MP��b��VA�gp"CQK�U�,C���x��M�5�_-��d���n�Q�]$A����J�����"PS�E���

��˸�.Rt{<V<�����i��x�W41N��M�[���QL�򁶴�*�Ie�*���eFF=�L�E����Qv?��3�N-><�f;��Q|�yr�S��଱�G�$�߬�33|����p�������0�^/O7�Z��$�d @��H���m!��K8&�j��_���o�S�O?Z.ɟ{�e�O�����8[(v�H��F�wT��%�(<ܺ��n8k��� ZzKÝ}Kfr�7A z)v9��}t��p�SXOס}C�j�{g�
���i����ג�E�pjo�/ ��͘ϓ������G�o_׉��u��>d��hdx/�p��}�p�Z��^�&`礓	�3�����3�C��pfOz�\�:ė�X���O�uu��a��EW�eP:���;��)ݦ��q�](�iiJ:}J���X��l����;Z<�܏q#���@�vY����0�`>,,�DՂ��V����F���+8[^W8�|v���u\�Q;��rH�?x��#	|K'�ӡ�`P�!A5u�ra�XYa�_��/D��[G�[f�D�Ops7�C�k�/			(ok�%˄�Ġ2(y*ݮ��d�,�@^�Yx�WY��:��I��Zm�6j��G��堑#� &Q��[�K��i.C���.C6&$h$��B]����l�����W��1�.�1w�g��ı���A�?ش��)8-b7'��>1bs�j���'�kP1=��	.�?f�rq��X����Y;�ȝ�a����5���#"�@�s:�;�<�4��)�ߨ9�n�!�J��Eậ��6"T�P;8�=.'`<3bI�` ���aP��e���������aQ@�AF���,��y2tr��p��[?�cEh��XQ�������VWA��zi����(����&S_�*�p�n�⊣��i�y���~��
2������$�J�%���L֩���<��0FBK��
A�O�I$Z�_0@���ő�<]*�h��Em�	���t�i<;#��,q��bv���f�&#HӋ0� �G�\�6����h3�|g��u~��L:����0/��W�ƍ��I `�,���}\s|M�l�l�t���4z{�'���qw2ś�R'�6l
����X5��NB^��䮒4��x�ap�$��b ���?NQb*$I��,��@."7'�Qy�zь\�m���-�����̭/�ꑥ�{�Wn�XM��O�0��������U!��j��F�>ܫ'����鍺FN-�ͭ2f�6M�k봾�[b�ѝ�WY����(�U�*�ju��?�R��*[�b^��8d��$%�Y3s���\��X""�'N��%8����x�w�{2�A{&	֙\���x�y7#N]����}�2ߺ!C�X�I��2����p��P'9� ��!H�/^;�,�2	#��+ǡIFo���� E'��?9f7K��z�B�dɎ���� 5lok�P��H��/T f|�t���qAH��0v�ʷj\]B%e��#�ѼH���^ԕ�'ށ��v!leW���D!TD��ɑ���"�g�/�O
��+o�mn~9[�PgzHIP��pm��%S7YZ�x�v��zI�)�+���.�:��)�
)w,�G�C�ֈ@bﮯe�n��ݣ�;��i^�B`Y6Jw�gfv�s֤�q�S��֓��4�ֱk�9�(wn��F�nh��,���A̎ϱ��Bx==a��/7FX𐭛����Nmx%�N��=5��_���-�m�|�1��Z���:9��?�9'n�ݓ��<aU!7�+�T��eV�h�c��9-(M�q �� �ic��|���{�X�Gj=��ʞ^��1�X�"����!�I&􆪽R-�+x��sU�}s�Qҥj�ֈD���$4m���d��Si��M̈��������}X0�e~UT}�F �G/����vP��so,D�Pc�3��"����
"��J����9�O�[Ef���rf�q0
;��#B����9ȁ9�HW��C�!��Ή�R�(t+puqj-z�	LgV�soU�a7B�X�����O��F7H�~�U'ԫ�:��^�F-S�Ꙩ3�6YA��T4ZT�]Z!�&�ڑܧ��33�\	�Qg$��B��@���F�q=��������cKH@�
����2�W�թ��fSޜ�9��PD��֝y�_�M��ݨh��յe����(��  �����(2+;P�<��4zj1�z�??~x|�oY	��i�P)��Ʀ$�F^
��ͺ����_vo�g:C���Z����J�h*	П�"M�F.����IG��ٴ'ت��j�R���-_A�{����ю)ݿe�5_m���q����c�l/�K��B�ˇ	F#�|�a�ı*b�M�M�:�IDn�W]��:�K>`���P��s�������2?�,���K'��f���/%:�Б^�])$Cg�;�>��`��.ZJS����F�q��t?�g��/�1������t���ϖ�P��`�v=w��;�`����\�4�ѧ�WVײрNAG�_���V�����V��dR8�~��G
�dEX5�ȋ��j;ĂT�,�,T���<aɇ�;!���R,�2�4E�%�rE�f޼9Q,���J�Db����ߓ*8�Z&�z>"t�g��71P�s��a�^�����������懓�D�!@�76xy<bֈpFݟ��
mJ�g���R
V�'��V��7!�mQh�=�@)]X:�Z{�w%m������N�ϼ���C<� _\���w��B_wL�Z�X�������oN���ˬ��^VD~*D��=�>--�K�<��N׸��EҺ����qoU��J7��_��K'����7���J��:�Ɲn�D�= ]*�@ߍ��c^��;:�h|x I�P�[�\�g1y��g�����f���*�˞�U���
�;S?!�.I�CB����KKSI��nyf0�p���ʌ��az����.�0�끡�@ML�؝�v���rg����-��i,_�P�=Xv�'P�!@?4�X!B�G(n��A^���ҿܙy��ng����!�k� w�d�,�T��}�'��7�V���!S�ރ��o�s��C X����p��b�Ҏo��d���MMM�___%��e)pU�u!��%ki���W��A������|��E���ꜧ�svla[}3zh~�+�ң�ru3������BՍ���!���m�;C'��H�wbX�,�*.$�9���LSv�X�FTN�jKHA�G��j�_4�;�q�\ķ�ܡ���VR�/p���~LQ���/���
�`�����F����W�I�]�a5|te���k�.����������|V�PӰ=F!�Nrv���7���e�`� Ԭ9d�$�T�5�S�.�9bB���#<���՜��Q&f��p�����Pr1����4��{��� ��g�D��h�/fY֝m=\�;>u�+�y?�3��j��]�oֶN-k� �	����(Z�DQ]jጽ�@���r���U�I��'R��Jn����V�.\�c /.��JdEit%�_�E�|Z��������Jb�|u�<��J=���G���^)���q;�n`~[�C�A܌�_��:�PI�i�8ǚW`�\da'�ot��^,P�֓���=��7tx�� ��S�����OF(zfJ�슡`��G/=&속��0��D�E��ѯ���b8!�$"J�KH�V)�--����R�B۹u'��Ssk�P�gga�U	�L�� �қ��k��ʅM	M�542.W����N	.1��V��3hIr@
S�ǅ.�h����72�'�v4%��pXi�H�7����E�Ļ�"�r�3�&<�����,;�kH6�mji�	��q(#`���I����%"��]�܎�a�u��-�仟$�u�ɞ�ZT��}nêH�M��@[�E�$(�44+|x�J�G&��-��"Hl�d�-��fy!Vj4L"���"�{؋v��;���^V���~���{�]����)� HT���q��1Z��f�UwVJvd8X�ю��'1Z~ 	d�Q
���I��.sb�߾��d�� ��*�Y�Jp�w+<PoV�
��U�W.6�kI�-���s"��$"�K���׀p��?^�����\����8U+Ž��y#�"���P�~0@�H��æn}j஋U�i�t�J�B����䠕�/f���|�TA3Ź@;E�0� �*p�l�Ӗ�܂P`����`E��eɒ�_eu���� %�F������AA� �A)P!���b&����B�Ȉ~{{K%�~1).*2�;����/�J�U� F�����W���[������?ʣ�0����d!�UT]2i��y�9���8�ݴgp��࿮sB�N�=k�VW�{	��v�̀d�'�K=f�9e��td	l�P��> j��d['G��I��Dee%!��Lp!�γO�[�<̾�H� ��eN��CW��ѣCm?2�?|wy���P	T���$h�����v,B(R�{���OP i��^���d
�"��p�Ix�>N"��`���M�M���ws��G��#K)�@�c �����/#�x�~�L]YG���$LcqVf��	g��~)�A�Ʋ�B�Ӌ��I�<�>Z���hP3qG¦#��ԛ�'Q��B�J�.c|Џg��R�F�|t�J��I%��_
�ʜ?��*�E;ֈd�x�y�:l�	Tp.0�i{#s�5p���A��� �T���nKҩ���╙��R��{hB�ba�4?�����r�0]��
n�f:�Ma�&��R-7�q\���,r�x��t���2��¦>���y���W��M}�H���h�$�9Z"��>G7_R�u�i���;��V'��[YF���nD�o|ň��O�~�����Ϙ�X��~�1�!�'P �E�K�ya ��Y�p�J����`�W�L�S������"�a�o��~���`�.kd��vo�ej���Բ!�.(Ŭ��DFux���@���R�@�o��??.�P¤<""�Z1-պ�ߒ�����]vfō#�o��Ȁ�a35la >j�WU���- �GiBf'vu_}�"��MW��V3������	cy#�¿�\�c>��#��˲�i*M:�c�,][, ��X�l����� i�x�*!���#U[[y|�����O.�&l8��^�aB�Z�����(�k-&,���U#��?$�uH�4��	�#��ҟ�Q�̬Y�4��0�b
N��bg��T���H�ˡӲ)��9П�����8sqج�D�I���Q!a���/m`�ר�Xe�p�c��l���²-��.ѧ+s)l�Z��G��ڨ�rV �^(���7e��c-� �xv��Hrr��Q�l��1��L�P·�L���/J��ؔ#W�*�R���?�C���C�����337`�����g�SL�s��?d�X\j�B��EѸ1�px�ݜ�bfh!�a�6�c�%R�j��O�Ka`hz��mr��re�Yq�*�ڰ��f��x9�\0��#؊()[��<QM7��� ^�(���U��/�Bx'��6��^:�8�Q�+��dGÝw�Xu }�*+����	E�?K���VPT�2��S��ȣ�&r �P*�(�Leik+e�R*_̝&���;��&��>�zA0��MWh�	�t�8��*��r$��G�$��Y0i�����ֺI�\�uXTa����.��R������Fi��.i���ɡ�$��l�s}�y����0��g�g����{F:N+�~���'�}j��iӢ��,S?խ�c�N�=�����Ҵ��K�k�Y��1�G�aҙ}��m};6�|�,y�дH�"y)4�����A�j(ᨀ�E	Q��ڳϢ��L���G2�`>Ç(��\ט�՞72���96���d���������Bk߬}_у�f���>d��"S?I�\����
r������p����kb���2P��ҊS��\ҭ2	���.��:�T,S�ꕧ�_���7�-� �Y��떬�kjꑨ�CU�i����B���x�}�����@�wwq��a#�C�k�O��>̕pUY+�-�%ӂM�J���}0�PZ ��ugv.����A���m=��ף�G��3sdS0��Om�x}��A5�*��Wk*��6k;�yT'��/�YF���Ğ������'�J���SJť�1�n���Q	]>?������+���9�e�Y�!Q���bо^��A�2p/n�~�2��j�s��Ǧ0�ܗ$c����O�U��hA���F�20����R]�^2JI�����l���'i|���H�m��j�\��yCC-\E�9�I_�nxw[�w�0ҒP�Ґr���*��>�mL 1,�!�ȿ����u�'	NGhy�^�8�e#�:�
�1n��a��������Bd�Dj���Z
�I�h�K���%����4���De��(�J-Ng���eI�Jj.����TD��-n��ieL�P��P_�7�[�ڵ�Y�}�I�A����L��V�(�S��b��ݦw���9��%���y���鷾�|��0��� �u	��d9	]��-襓n�� QAl"=����%�cu�c�����^;u�^��$[�"�_��&����0��2��;���>8�;�؜�ێ�c}�b؍�&�;���6�8�!iG�lhL�A��:q6(g�.�@]��s�$�ee��ߔ_I$@���B�m3֔5q�{^;��t*�@��H��
QI\�����l��d���Y�uL�"Q��I��ޱ�u�)kCZ0��(��K��\ӏBŗ�%^B��H+�w���*'�n$�:�Nk�)D�V�r�,�~jת:5�%���AN��P���Q����� ���ɥ�z�+uKC��D�BFJao�tڍ�:Ӌ�)3��cL��!���|�x? �������Fd�<���HZ���Ph����v#bQ_,d��o� �2�*$ �jx�S�3g-Xa�:e�L�̅e�;$�,�o�O_K �XU�]&�QY��_�$td��Y�2���}i77o�}_�$[���`!����������7o�KtB^ŋ�Sۛ��o�J�c��U[�YB�m�̦{<nL�c�8��l)�w�#V{��!Tl"@�V��M�TD

�����^ o<�� =+	�4U&��ż��?�r��E>��Oύp��@bW/�) d�k����t����Q���cl�Y���D)YX)���*�C,�t[1�d�\�q�ک9?t�?i�q+�y�+�=��8��t�=T,�7D�)lX�')Oʰ���a�W����z}uv6B��j�M��rRE�W/�Z�����Lζ$�-����S����ү[ߠ�^��k�*^�ꔹ��L3�J�>N�,o�H�&[�)>�����$M[{{�f�8�y�6z����3T�|� ;��ZLl���œ�Q���M���_��g�w� ���W:'�o Ԕi��"��)�h��r�{xDRC�i>�w6��������!>�u<3���v_���u���ص�4E/g>����x�6�[�G�K��5���=`�dfvd���şy}*in.���/�o��̈��D]s���ד�'�2Uڅ%%Lud	g�ӆ^�����
�E�dt]oة��烖��٘�I:U^�-kK�|�	�pȎ��"���^�QSx��$^v<�Z�~Lr��i�J�GvL��|]����$�REw�͑�<�sӦ�U��"���G�KT"&�L����}?2�hR2�����)��(-�Q%�t6W�$�8I�EgI}g۸�Q���c�q�$�K�p6��?�Y<=9�݂�D�IU��xb!���� �#n�Y��ض'���C�&2���E�<��O�~":��7q�	/|O�s{�陯N�J,�>c��#��E�5�/�q;KP�l*�b�-	>�;ZH`��_lΦA��.*�j�@�*�ia_l��m����n�(�*�{	�v*�($D۸��9Z���'�?G�7�n�WuW�K+� ��X��i6�����1�A����T��J��NZ�����S,n}t凣��-{��\�v���}���_O�uĜ�\�|� ����Su���kWb@̛��9�>
��P����:����j��{�����7?���_��*����*��F�%'�K<��(���:���a+���&��4 �������0��긎4��z����o��/�]�ގ�7���E	
�N憜��0��S9�%o�S�������	�K��wv��d0�1+8�3c�6��x9�m����h
�	篷���������$D�(���K]ҏ�����I?j���p��w�n�	r��I����d��Z1�/�C���E!��q��OY�yQG4�D�Њ��E;�_��q��ba�V8X儐�7�L����=F5�x���¤�ͬ�B1>z�i��[�xt�&Ȧ��+;��'���� ��v���\D�$.��Ќ[7�;�u�У�A�_�2|�o	��^���w�/yџ1���G�a��~��Z�K�	����,�A��U��Z4�P�By���85�2�%�^Wl
�l�ǰ�H����Uc�Aa����ߋ�ta�DFf�Ϳ)_�i���z�����������}��g9�����A��US@;Y2E�OE��k�s��hrU�Y���/�8��L�k��D>�|su�@�i��&'U�"=Y�Z~��+���u���0p���|V�<+�l(�4R=~oVI�����b%�OI�H
\��^�.6fnj��po<��L&2+�2*BXI�������J��˸����a�W��V���-�t���gB!���k�;:���OPǛ��]����/ȣc	H � �ׅb�,�I[��K�ԓ�B�BfN�T��$�j
�xR�ƅ��̦���e�#A2I(���z�Z���LQ�����0n�f�V���k�I3�DJiu�5�>ʩ:C�T\eG�J&��롻�:=l���!�<6HzԦ��w�����"���ؙ���[+��4�?.�v)w�y��E�e����Z2���d��e�N�¾�?I���&�@�9[��H�N��"�m<L���r�� [�y�A���[ДM4�ϭ<(鉸���:9T� �t̜�����-N��6��/Bn\t�:W����_��O>����T�P��F���|pr�2h���q������:8|R)��)_���߸�����f���g ��׶���r�y�v���ɑ���(/b���C!����%���g���ө�I�yU"v��-��zwۋ��y�2�!̦��}.��2B+�������(a�z�����P. o��<�7�/�zE|*)E�H��%X�@�n� V��hs���B�ꁚ;��Ǿ���7Qx]�b&�F{v3��Ȗ�0 ^��@�����Km�� +/�,��?���z�~\C}����K$��D
-�2�Gt��!.~t��CjX�^��!j�( �f]X;*���)LH��#É�d���Pv8�v�y����������Wȿ��\�[�7gϚVJ1�VI�����������]�X�o��YA�X�
�q�5��
n ��!����8u�x-y�{��w��Z�~e�2�ɴ���z��Ee���$�腧��N1���np`&!)���-�@�Bn�Jq��~�VE����w��Ǹ��ӿ�?^QkX�Y�>:�;���\J��
l=��-:l��C\0������{�y�����n�q��\���*��S��׋���/2��8�:QIA�1��D4�4&J��Lm3��d�p�7�a9�a�_�;!��L��p���a�aw�
�I��6�_��[�-1�|S�2.vV���+����
��p9����z߳1!Nɕ�PG�v���HkqY�n�D.L%�ŸrO}� ؏���Po��e�	�(���� �{�Gԅ����f��"��dy-�\~�DM�<��_e.�}׺��	o��ҫ�U�v�(]��1���Gm�`�f�����p[��"�m�k�_���vw6B��|*��6��z��iA��Yi+(BGR��� X_��Zf?5�8���^m9ItN#�S�o�eH-����.�xr� Oa���'������a�,�mhD�]3\-M�6��b4TPv�CǫC+>O�%;1�����S<�+$䗔H�D���5F�V��蛊���~;ݿ�Nd�H���*~��0~phQ`{���`���gۤQ�6H)�|�(���,�(g������Y�Ҫ_�՞�0�$Ĩ�!C�>֡ ��v�I�/�Q�q�����j�����>����ggO�h2��������daй�`g���w�MbᜌX�q�)�ʁ�5*r����Z2�k��K�����:�_�QNE��H%Z�r��0J�Y�y����`��^�g�D�#3I��l��]�ݻ�C��p>��,�}A�N1��@b�[�)�N�|���_�hDu�������$��ӖtM�E��;����%�{U�XX���e�2K岫�K'Qv�1_�ε��yh]���(��L����r�<��iΝ�i���7GdI\����*_��i6{3&-5=e��t������Ŏ���R�gen0���.����3��$���7<t�z�>E�=%˸�ހV
�=y~�"WpAW�yT@�͋ 4�_c^%$y������������m�A��'{1�������h��60&h�-��,RL?����w���$'D�2����p^����5kC�Y��E���|pު��5.'˓A�8 4|�&61�M!%(�'d�ɾh�|���C%z"�gw��?��!�I)P0�ɔ�g~<6�Ũli���zn����Fu�ߊ���%��EV"��/R�xK����?ж�y!���@�[�|�������z�2�a�Q���bs\eOnj���`@	�O!`�]7���޽܈p��u��)�;�����P�7� <Cq҉YZ����]������悸4����ߊ�&��1{
�c�I1
3�-G��-�~^��A]6��: i�q���'�^���)��W[RI��H5���q9Z%�=sY}�E��Z���+�P\Ȟ�hoS؊�D����]��WKPOl�p f.})4�A 㴕I�c�r������ؾ �1�׵� �#���%��LaҞ�y ��QR��� �)j����]B���*��u���FJ�\>e�p(�n�����CD��Qjѱ��w�
a&s�Z|i#n��]o�"1�)6	i����`S���~������o���������WhJ��e82���b&T��C��E��N�v㧌�:��oM�[�u%����E9+Q��"tδXTUt�9,�g���]�������=m���2�-����pN�o�p�_���9��\% �-{���.u�\<{~���F{LL�"�ܬ��,e��2�������S-��rk�o���lLɨ�{��p� �����pb�v�5���u��s��?㸫6I��J����t���x����<�+��d��n<�ôy�N&A��(z/���i!�@ߺ<+��h�aѬ�MX[���K.N��6�X�XhYO��"����=�;#����-՜_��t�����'�!���r�ʇB���"�h4s�Y&kk~5�0O�D�8��A^yy!Ȣ�I&��^]F�0lY�{��Q�j���	$��<'����=9֍�11̺j�$ܙuD@hWC۵5w4��1�q%�.�~�qD�ssٲ7?�.V�M[5B��d���-��}.!|��{��I9Em`�,���7/�Հf�>���V�ņ�+���7h	���/e��(����O"3��I[��]�E�RU}�ʁc�x�J�r��

�^�
�e��t&6��L�o}%W�#�9�����X����E���#���z�kA�����x9G_")����YBz$ӝ2G�/j>Y(�e(r�j�D`QL.�ƹ�l���4��Of[v���T��iߚ���S�<.f���>��Pb�>Fb".�?pb��j3	��{8+@���ТO$�Ύu!ϒ�"nf�� $c�ܠ��q���L�:��6R�꿇hX5k��6�Yn������Bg����{����>���`U-����7K������N��GB�������.��̾=5��-�����?���@�����'������N}��'��h��/�����v�c��X��U����q����I�����~z���;��v�\ig��"�=[��ޫ����0O��/:����l�O�+nť��?��Uj��>z 7��-����P��U��Ԃy�*������1�Nz��Y��Y.���e�8��TW������#�(�6+Uz�+��c���	<:���խ�qs7��o�ֲ�o�����s���V����&��p�ўֆM�1��A���qƼw~����'vB�_|�q��MeF��;��S�;4D��޼2���ݳ^�ʎ������������T�g�����iUGC�I��f�����ßt�X�"6t�h�4�x���}A�U�		o�F *TR�U�	t�������v��1�7$0CkL�6
� �� <�tzF�op�2:�Ъ� f��c��A�V�~���s/�C��+��#V(v`w��r3�]�H�p�Q����f]�!�ݑS��B��+�����R�۵X7.w���`��܀�LD����ǵl,�)���e�4�;@����Z
�_ѳ9l,e���D�m@�J�؄���v�5C$?��	����q���7�J�lË�����G�q�ʐ̑�ҡi���D5���m�s�!����� ��ĳV��x.��Ӂ����*Tz����zP��Gq���q��ԅB�v�`U�MUY���F�O������`G�xY��MX?�`����o�RF�Y3�r:�\	��hA888c��Jׯݦ@�i4i6�kꗐ=����O)���s��/�4'�)�bY��t��r����擡�9��KK� 6��ݓ=�&#�+�{;8����Ms�������@X{�ЃD {\��;�YO������/be��*�8�k狄�t��t�m�ː��t��&�}9�ݱ5Jj$&�rb�L�x3.n���X����E"��a��2A������+;��yg	>���_�e�h@gre��[����w��(���m{M�<�F�F'57H)��3��D\h&��Q�(YoM�ݯt�b"�������L�_ ���p�_��k!�����Hn*k|d�6�g�/(e�Ao��>�=;:���m�����x8�>��$^n�L�mK�e��|�ܺ/�C� Fkc޻~��;W���~���]�����M�����y����d?(j�;��9Gdc��,�;�ꌃ����S��oG�;���	J�gư����<�����V�����x�rr��~��HE��a�$��l�hi���d-�ը���O�'��r/�~^�]�e޳�)Z�_	|U>q�%l�߰�<")�|g�H��k%�>>V�F��pq����Llf�J`u���Zo�	m�3.�n[�4�+Y3DO�V��T��5/=��ϓC�����|�&��:b�jgr���r.%/hVt���NFF����*j�U����G��������x��;��(x%�f��������~��$,d*�x��]��~C���yj����Q���d˭��Ź��M�J�S��4�����V񏙥���F��6�Lc%�<�~��+��j��-Q����=
t�8$��@�}j|��r���;Ў>I��ն��or�;�B�AS����V��Ws���4Hοt�zk��E3#����~i#0�<��'�&�V#���^��g˻7�SP��Xƿ���c�=���}������/���S9M�+��9��z݅,,���W ��O�]L�L!��r�-(�MV멆�<B"w��z?�p�<�u����R�MZ]a���wd?�%{\��'OIK{���zr�ж8{�Ѕ�ļ�Ź2J{�7�N�U��^}Nc;�ypb�T-ZYu.OGL����-e�x�h�U�])�!��$�.��c�̩�r>�[��b���7�PJRQ��j�_?��5�'B�w�0�=���Ɏ ;���Y�O��؈�&��H,��-I����j0�&��C#��D���=�-��c�����MhH\IA-�xqj�P����J�����*c4����m/]	(�@1ZP���p38'Q}���-�8�=����ԯa���ּ�����^ �}3��\�/��N���U"Ρ�1����t�k킀���C
 \�ń�d�:��2�]r��V��.`��`��eyGZK��S�f��+�f�ٮNo,����X.W)rs�ʒqҘ�˭���Td�,B&�6ǠXf�޾H�� dZ�����5QG��1x�)r�k�'�K+�Z-(@<�{]Ѩ/FI���ho_�k�Rm?�o���Xծ�~����>^z�5��sr2��z�Z�q333��k�޽�[�>���۩�8zox�x�u�7����&X���@Т�����R=ĕ��]wr����s�u����x���da�V"��#G��cs07��Սm���c��P{澅�����
	I��&��{Ʀ��p�i
%q?��<'��Yr����Ȣ�Ǹ�4�~v��^���e.���E��Ѳ^1�3h�k6��墂GK;h`��JfŬ/Uc��9�4'i��V.�J�X�6��8���)o����y��uT���h�?7�-[q��#��fz���	]]����|�(i������]:��=�(i�6����,����i��4����1a.����>4����z���Q�*���4r����k���Í�ed�{?"�h9s��CK�A �.��uI:;,��ꨏGRoT�e�i��9�ݠH�'�m��ŕ0:pO}w�{ܭ�.LJ}>d�V�o!Mlgh\jM(�]��nX齕N�0[+�yă�}��	v1��`ݕ�R�{�=����xJ]�[5�Yɜ�iI#��Z�������F���<��q�ը�;�E���9�@�`��V��0M��_��!�D,i~�.�ϓ�!�|6@�GT.�s����>��fA(����k�;����v�@����JROѕ	H��/O�<2A�N���}��}+��rs�y�����LB2����T^w�Ec�N���nb룩&^_-ƞؔ)�Q�{R.�6�[Y���u�Vp<�j.tq�Tj�tv�"h���a�A~/�$�.�0�{-9�Dd��k9Φ'����j9o�El�����-�L�Xz(�uq�?K��hv����%��08���+��l�����������=���J���K��f]q�[]~��+��$j}�9��\]�l���BGv�D���eu+Y�s�wt�~�(���{��x`q�8�B�r����R����0�]�C��p{i��BF5Q���@�+Ɖ(4��*`����PO��wu����g�U�%�ܧ����Q���H����*Y�r9O�r����{7�Q�r	C7X��4+M"����g���'���3O���I�(�}�#z���#z�Ǳ�i��sa�%��B>��gm{��^V.�G�y~-�뿠`�'q�MN:��,94\xS%�Ԏ�{�HzX�=�Z!\�X�T|@ք$�-�T"AңQuow�t��ݤy������c��X����]��ūˤϲ�[�/��s�ߟ���^�9���Q��0�p��	��)Z�0Z[ܿ6<2ӄ��=xg��aP����K�Q��̩gt����b��R�O�8�_S��\�ws��6 A�h�p�{�En�7(4�BI�]�B���uPq�1�k[f^�{>i��7[���1���Ԝ����9��`��ґ}&-݅+���S�z,x+�Y�~(��ku�t��j�~�xK���G�qd�z��{������}�� 7�����Wj��rD�sp͝#�z����O���ʉ(�8I5�VIr����7A��JC��x�vyՕ�Z!��H�,�̰s���r�������8O9"X��f�[����[A�����;5{����fn$�eR\t�_e��*}=�0�m���z;��0�B?kDQ���3l��f��h�-�7��]:,?��� �D6/I4�G�D��V���*YYS�e��I�@���M5��o��k��ty�X���D5Z1� �즊��E0K��p 7K�b͸R���� )ᗽ0��Ű����u����'�>�$Xꃓt�j�iaQ"���E�>�{��3+�7���X�y�i'c��[�m���q�d��^�-��:0�9�$�l=�b�m�?1�b�iq��f�O��s2%]�fWv�j
��-N�vF�|YH<�C�t��+����ֺ �ė����c�S#ց�����/���yp9P�QP�l�t�>[
F��z�\�I��t��v"�8�ν�BV����5	���\5�v�=!�MLy�8���V<�*�_�����h��Q�^���f��Ǻ�੉+r�_
��4������q�zS�>Ï*�"`���"H��	mm�6���ԑ*�|���B޿Q0u(G|�(2�JA�*�w�p[�u��sh����V�	��<zW1J#��y����#��fXmcOWK_:^��LO>�נw���Z�x�����ԷZ��gSX���à+j�d�{�Q���p����Rk���$������46|��'Q~�ݫ��˓�\ҷ��pP�PX�v,��^F/��6!1�`�^����0Ӱ�&A'N�S����`��8����u���j�)n���sT1�c|VI�&�={.ɟ��z�H6�5�D�%�?�/|x�y/t���2�J���`)�����:2�ސM$����ã�k��h�;��o'��bD�H�:��xY��9^�CrF��"C���m\��\a������T����zؠ�ɍ\��K�n:��� �j?��4��b������oJ�6��Rrq�9��d�8A�vu�C��Rg೩M�F�á����N�J8��߰xK�~��p)c5<�ϟ���4�* "�D�6�([�;�s���v���Ft��������F�>@�`��p�;��z?��<�U'�����{������3j���_�Ҍ�<��_Bc�\�~�cV�bk/>A|���R2��u��D:�uYbd�t'�W5�~��C�C����"z�X����@��3��6�s�l�yg�.uq!f�^Y�I8�e	��g5�:]Ȼ�T�+,�{����/���Cn��Z�
&�#}s�����k
ȓ�%0���r�4DX$�����s�	F�8\Q�>~��|h,ꚳ�8Q\ϻV�xW-yލdo	��)�W;!��郛!'0?!�O&v����j�9�����*{<ثV��*�/4���U�%q����i�b�l��d�M�i6����TT����.{��>����,L��|�Hr���%���!�{e���)3u�_�՚W�F��9��z!c1ӕCv�c�Q^ћ�O���
�2���*�Tw�HZv9��C�}��)퇞f����e�=>`��56���;G����JV�eR�|�?�p��u�l����j���&�U4�Z#�����B��.6��c32ti��{�a�i}�����K��0l�[�H�uZjk�f��[)�DO+%j�Qy(���_C�����W5\�-�5�d���7��|��ﲇ`f��f�$��!�(��P@>!.���M^����S�7�K�͢K!��庰=� �eu'���~�]�J8�P�If����EKy��[^�|[~�B�{��SC������t�w]3�< ����9�Z��?\-�B�n��rz��U�?��1Q��XfE��h0C$�Ɖ�ƒ0�� �P6���뛄в��ߙY����J.�D�L��*����(��%���U�d�l�q�̵�q|ϕ�zT�����J�LE�5$[m1�7K*21�=���tƎxb�\Hp�t �l�>�L�ç-����1���������z��e���s$Ił�ǒS���]j&����;ҽ�4������Z�������9���������H�$l8�i�� �L��O�=?��6m)�8�XQ�y�-���5���S��2�ˇ뒶H�̇��������䞷�.���i
��;�/��~ ��~��$ٮ��*H�W��E=���ڣA������K١�ͻ�u�.Uy�\�<��WK�+�.�F>�7�җ���>�c#�$�%�ݼC� �.n[��^�m8X��q�iG��0[ȿc!�#���`��-!xr�����rt��X��>��	pHyr�ڙKБ� Ž��f��@^Ɯ����v��_5�;�wg���<�Ȇ�a�O5]�n�y��c���W�٪�>ɷ�
5�u�5�#_U����ʪ�'�Z�n�����U����<L���V�O5����L���{O�<Z.#Vl,� ���Q�?�iВ�y�^�d��Kˢ`&���t��`n��n�jz祦�m�����KPQ��m���T�A��c�j�A�첿/��US�O�KO���S�w��V�-�dBl���7/c+j7��ʅ��z��xu��[��A����B���Cu���Z^�yHҜ/n*��y3�|�A5�\q����{��HN�.����L�E��8P?�hzZᗭW̌lq��:�ܪ+�G#���Ê&r��ړ_2&�f@�|Vw�4G�I��py����v�Խ�`�8�[MId7��p����:�'���(9�^a*t{-�B�22p���a� _Ym�m40�S���|h9䶮U6DLԹ6�#�L�RJ9z�`��d`��91y5�,����wm2"p�# a����j:v|�s��B.<)#{��pq
f��7����R�H*�Z����R:�'W�#���é�!N�ܔ�gPZ��������S��f���;� TUh���vL�|gB�}�����3�ǂ"��� �57$�oG��1�a�!F�x%���7�'��Q��''C�U(I=�򠉨���Y��@���8nu+� I���Y����{�;�Y��0�/Jˏ���Ҵr�N�j��'�ZE�ߐ�W��=O�p�i#Ks�SQ��Hݵ�t?n�2����츙�ȃ���>�چ+ݴ��r(^��xQ�WW��FH
�d��C�c��+�]?�Vjȷ�=c��A�'�HG8�K�'+����cK%�J�@臐Y?��IsYso|�̗6�K�8aT�c��|��@���Ǭ}����N��&.]�z�L�|3��L|�x�j�����ٶW_�� \�r'6���k%�=���\�[���g��S4O�W�Q\r�(&9n���J�ux��U��X�kMm���.Z3� �� q��e�#p��j�J��<f�W_��j��C�l��(i����O����d��&ЍU�J��u6�g��+P환i&�;��rJ:ncј:����u"#�M�,�����E���`.c�� I�WM���0�n�'�c,K)��]%)�i�Ԃ&�ʩ�����IƔ�pR��OH�E�OS���^}�F"8�(2Zyc�`��q��x	$����1�����3a�k��c �G"���W�K�x������$��C�GOĽ�9��ұ� {[�_��=[|@��:�h�~>^����0�|-�/X�����qV��z��K홻��R��$�i#��3,����EH������L.*ĥY(f�rp�)���9�7�]��@
���O˻��>�Xʋl�B�Ŧ�(�j�Q��[k4��)�͇W��ݾU����x,�Y~+c�+�T쳝�b(�qQ�N�GC4�5�^}l��]��ѭ��yzx:/�v������8���V�@�<hsza����!���B�K�6�(�dQ����G8�l��ř�a�A�R!��c�V�]5����F[��l|��kKg�T���jR��hb�o��V�U$�0���@�Q�C"œW�N��_}��vj�� �.?�`�:�sWvY?	�D��~��Z�o��<՜Ay���N�q�~�mo��Wx�~���CQ\h�N��ŕ�)�������/<*�:<��5��C���8:S�g#ǎ��>��@�zo�$f�|=���;'[�����->���w�yBi�'�*C��%e'rXiN,�:SV�R;�Y�%��xE�� �����ީ�[G_�Z��ҷR����6J�E��SԵ��+�_��ǢJ�%^ink0z���٧���\�DU�+�K��G�Ѷ����tO1��'��>}�&����Ȼ�/	�����c�=ߝ��K-���ٿ�8;����4le��Bf�'��L$�����@Ȟ�O����Ec��ƀ�q�a"�fX���4�7K3�>��VH�tY�%�߫�?_�� ��_`A��4��ӱ����_��y��R8.j�Yw��vD^6Z/�a����Ɔ(����Ęe��J��$��(�%?_�G�H� ��q��k���,��;U�ˣ��J�B����0Z>�L�rzXπ�%�in�e��Ǐ+���׹�V!���aB�[M�_���������C��������靷��k3��d0��<�\ԏfVy!�b�h��ln���y=�E�����XP���XzX�%��C~l�;�ϡ�8�s�+��6s.M�8�*�������M�b��x��:�����v0/�.$ҧ8�_���E�����TL��m�~�*B]sf;������3�p�2��V�b2Dj������~��XqIn�j���	����}��l?03�t�"���_SL�7��"���	�?O�Sy��W�1횝.����,���b�m9#���_��\�@�6=�'ƒ�[҅�^�dm��Սe�|���s!/�׋jΔx��g�WzoK��HY^���V�{�䈉ʑ��@%�G����"�"�Isp�y>�q��
j(��������v��� ;y��@���ͪ/?�ܙ�1�W���y��!�q"�(� ���>X���s�'.��/󪸺�
W���H���T��C#�۾hLG��K�xO�C�˶l�h*��wwj�g�t�������5�������԰y�螔5J������!ɸs�5��#��KY�VU�I��߻u�8Qf�|-@b�o��'Z����+3P߽�:�� '�Q�	��kh� ��A���57�CE�׸Y����y���4y�	 �QS�}_��.��ɋ���PR�KO���Z���:_bm�EU7bm���$w�7K�sX���^�/���^�'_���nwL�^�G�E��ѷ{r	4g=aS|K*/���ؓ����0��� �#�*�N}qc�oX
n�RO:�ܱo:��mjN�J;=pW Qv9R8�;�5LRp��0l��fU���%�L
S#��YL�g{5�g�yB[=�װ�#r����q�,8>�`ebT|Y��u��gӲ7��?<BͦNܵ��{���RA�2;����1��vc�K���=eŞ~��.	e��b�����X\9�ߣ�{FU����N[���m��Jo"�8o�ޓWg�!Q���ۼ�zb|S�.W�=�ʂ�Z�H<��uk4=��Á����`�Q-%��}J_�v^��\R䢱��3H �]�����Ԓ�p~��АR��ld����N�`�(Uj��d́c���#���۬��,���S1N���农u����^�FC���;����}�9W�?��-�J�e�%�<궄�7�c��PAөo��E��/�N�<.ڮ�A(�.Z�Мr�Tx�N]'p���!`���N��5I���R��(@�Am\~Y��{�?��;����j��:E�z����"ɯ�Pci~��ػ�����E�5�.�+�$)�)����B���SH��o	d�i�N�R.D�%�	�U�e�Ӈz�慤��_(�J]��R��:ՠK�}z�P�����:�� )�(�1�f�.DU-h�jj��K��	Qf�Vcw�n���4��,�2��k��?��Z���B���V
Xc7w�b�g���"���.6�ˁ��L���D�Te	��yY�8�x٠��>N��{~�N�'N��������,hb����Eb�ZVFywPMR���YS��9i�5�y��C�l�%�	���(����MUA�D:IIM(P�Vl�[����$��;�ZZ�)���)�eQ��b�okU����[Nݸz.�q=M�_=	���6�C�Pvm{�HZP��������/\)Q�2#SZ�y�F����:��ny{�ҍ )�"]R"ݝ�tI�4HIK�twæE�.�ͦ�$6�����w]�p�Z3���Y�&��� ��ƚ�y�ޚ꙱M���>�o��UWzY/�8��+�����@&�d|w+:7L%����#�ؕ�݁^
��|Z+������犙8��E"Ƅٚ�a�4�#//y.��)lӦ��)�{NO3��j�)q�U
��:����@2�wǡJKl+*v���������8��2�!B�s���[ W�c[�#Ri�T_���!r�0(�F��3{U�\E���� ׄ���9
Ĵn�9����������[k�q(�č@��o�uI�m�ؙ�Ւ�j��P9����MAӏ�A��%�$!�x�����`�ѐ������s�n7ov�7���j�t$s��F���h���{��YdD�wa�A'�l9Lh٭eԽ�O����0�>R�s�d��%�C�����T~S%��l����-�� %i
@Ak���ݼ!��jb��U^)k�l�t/��*k%nl/x�LD��Ш��Rp�׿X*Y��(�a{y���CU�.�_ٮ~�БΕ�������i�b�?�ޏ;��9E�\�`t\W��juH��X�4̴?�zM��- �]m��2$�e��ܮ���ދr{�c	,�'|��0 �/x4kV��'!9>x�0�BmBj���m��wSGW?wx�/�6;Rn:	�T }�2�r6F]|��)��=iѓ�м,^� �2�ekr����;!�t]@��W���W�	[>���z�|ȇ�\X�b�y�W*��Q�?��q^��%-y��\\��ÝK�9�g7�?������2,�-#5�Z�B�8���Q�ůij�iz�+QϷ�׸�R�g}{��E��Zm+s��7��`��(O쾡��疒4�7=\n��� ����/�uH�h��hli��3VEgttS��A��m���._����n.�+fc��s�4�?^8.O���6̂|U~d���{��D��o7}�E������H����ؐl��r"g:I"�`f�q�~k5����R*���I
���������"��q�LZ2��������g��<,H�1rXw��U�k�')��4��k���\�5l:;!&��8�4l4$.h8@��&��|�X��A���ƽ+ᴇsn��J��ae�����E��$x=���T��3W�ش�J�.	�h�����+Fs�	���\jL[���Uuf���_ܝD��|�0@*��*��qJ9����$��W���'�7�6W���?Fqu'(�{�D/#U�60��������7@�ac �j4yb��>�BQK8���uA��C�QA���$���-E�
�ar�
�-h�AILg}��hn�3��&Õ��, N/�i�0S�_o�7MF��К��n�#�P1��Vۄ�O�?�9�p(�����מ�7Cpe<{���B�tσ,��e*�����������yM5���ƥ3	M�����\I��, /�o��a�qBVtР�J�k���i���
���r����ϯW����&�-�K�Q�h��K�׶�Z������A5G9��.��`��}���]�,6��X;�Z�"\=}wV4�݂?�YR�Ic�R�9��z@����u~���+�hr{��3�$�Hb�w��$��3Q$��q[���8���_U7��V�9�ck?�O�����lo�l����I�[a! N���2�H�?����|]�f�z�gO��Fg�!������W��B.���2����KT?ˇ�:��d�T#J�zi/d|��Ղ�:���6p^:�s��:��ٟ��M �tCC_F��/b>'Lb�Y����=�0�A��F�ո��qH��jh6uF� ��=�X���8xX=bHU�Y0VD
)�k~�~s��SSR^��o'v��>m�HD,U�(sdu�W@�������P��_���!
�a��5)E�Ӥm��&I"C��yg����`��=p�n�er:�����0����)��ܐ��7A�0D��:��W�\Յ�|�o�e,u�s���[�.��u��"�1�h�/���yd�#��45'(������@!X*M&Z�l22{/��Fɔl<�zZqщy��5�*Qb�R���B�֠n���-�xG�a�G�\(j��ȼMB`t��1�)j�0#��{��͌�8!ms���T���b�8M��f��0�d%fDg��e�$��盀�Ŗ�"���!�?�W*�Jc"襠?��Ҟ5�8�n�#���� m8ؓ�����-5+K�R�l�c�x�;�oו���g?ONf�&�\��ג��a����B�̚s s�%	�|�d�z����dlhTU�x{3V~�@8�]oU�J�4��&S�?5�L�;C�\,'�
�o9�y�o�_���%����{R�'M�Ϳ;�"���9I0qQ�W������?�~�=Xz�:��$��	�J����K���M�	�s�!�S����履�U�_H+��L���f�*�B!R-й�QE������F[�<��\��*��9���JF��h|�̉q�3�<��qG�n��)�Ŝz�k�M��/|�B+�+|x4_a)j�����~@�r ���Ŏ�x�ST�~WZZ4l�x���$$�H؛COLMM�N�8��g��&H����i�s��;��Z�}�Hɿ[���D�x��7�� ���Q%��A�5��j��cJ,Occ��z�w-�]�_&��kB�GK����=)�F���}�0�P�P/��T���)��k��c��!�
�P��a٢��{�-9��T�;� ��^����P�r�y����b�N��4cç�p��-	q�:)r�G�k�Uf!?�����o?x��Q���}�0
D<b�ǒ�����<z8PҲ��{�MZ�}���Ϥ�=-�<xի��hmBh�c�d������!ٍ�%d	6�Տ��f�H��՗�_C9�Aþ����6�����U>>b��U�{}��d�GH�7@qS>�/`�455���2~OX�69�C�Ar�����3�������������I��K"q8[o��W���5F���#T��Xw81���#0�{9/K���k��D	���|�ʇ�VZ.�E�y#��b���B�S�H>4��`��؅���ZgH0l�mH����M��!�.IN�L��?`������j�V���9Y
�r$u�����-|���p�&��'��;� �E��IyoOP��mZA����6\�m(=�.�R<Io%5i\H��J�������z��P��'\�� �/BLX��ZW�O.}>���u�Y X^�V�5�E�~+��߀��06�J:6\ܳf���2{z�����L��5�͕9��<RG!�5?.�Q�#��O��1��S>5=e9p˰I,Fan1}|�]��;&²H>^mώ�#��j*�Z[����n��֘�y���&+���$��#�窙\��@c�v�'E�	�����Zɧ����PM6��%�;��@ʶl�#�.1�*�.� �tĬ !�O}��5+�ԃ��ݍ��jꌌ/r�%T�4?dy]%�}_˛췪
��Q|�q�9 ��%�B �T[SNc���)Y�Ac)��J�*\��\l�8�b��D�X���x�k��gr�W�E�'l�����:��A��vՂnJԧ^c9y9]e��[���{��D���C�)��~��|���.���uՙ7��l��.�.�:��o'5K����(�ſ`��Ch�TH��r,B(LS���"!ܮ��¿'&fr,��Q�;2b)�E����F�o�����N\}�o���͵�>z
��֦����:k����UY�֢8�	>�e�P�"�p�7�E��S�}��$�0��M"��/��(���^�'D#M���d��7׃��j�l6OMt����Pl��6�����ylW�����7 ��:�Ի�������B��y�۔N�#��f���Ͼ({˦%C�� �~�|��!r����y����L {��(&`-�s���y��͑G�,)���߿!�h��Rb�U���<)g��S�hUuʃ�wvR#'�+}#x�<�{��w+#��1�y�s�Ub>��>�	�]�N��G��8D�j�á�J�o	O�d�U��im����44����'=���,�I����ƃ^��t)X sD�)�⏐g��HI�"�>�� ����@�������˘YcO�F�4�\���	���c�1����c�V���OWMƕOK���8�z���}E��"�aDH�!���!�!
ˍ}���G��8 �i�ۛzH
��<��K���ɝ�ú���͗Q>z���$�?�����3�S�7�����0͛���c��;��%��S��e��1�O�J��w�M��#M)^�1�{
�A^�8_^[��������>Ϝp�z��qu<�g��o�l+�^_�˕�&�S�|�2oT��9��c���k�E����1��������l@$#�~J
�*ɩ/>�m�PT��h�BZ>媿k���=�L��Ɣz�9Nz �z��iU�H������5h��m�~��{U�\���,�|,M�X�i�c��������j'�\�_2χcJ�?^[�d��K1�f� �@���^_��u���Gf�$��OR*ΑgLόW���K�}v�������@===s���z�a谆i����" k��
�u�z���Q$1f���-L��R�B���zF������BHc�=��fрl7e�mL�x�徝�`F;�� z�{�ž�G�X��҂D�O�ʍʬ�7s�eo�	������u�]k[c>r� X�`��Q��xE��T�,P"�F-prN�p�6�H�Jf�ցD&�:R���H�8�N���m<��'�͚ ��8̾�B�K�W���ع^�&�:��0I!�sm�Z�������@� �P��e��g�d���/Kewt�����Ǉ^!�
)W6�hj�d��*�>�x����ELf�f�w�:_�<1�����ʃO�??��?WZ�q�0Ӣ�:�"���o�����l/��4�b	���1pz+�������9��J?	�{�V��%h�a_.[Sν�O�	ܣ~߯��l�csqu��r�Sa8*@V_���\���=�7
��}�DR(�
_{��s��bUja�+"�j,�����Y�L��������l��Ћ�av�8�`W����pw���D����D��3Z:��@ՠv7��I1P��S����Z��:[ۼ)z�;�ڀ�#Cf	J���-����v�Ԁ8OO�*2j, ��e�����M�ҭU9��n0Z�jTB6��$&4��EjؗOgM5ҟ��Df�V�Qx��O�+|�	qХ�$9��?�$��D{s�M��D �C���oeޟͱ!���>N9T���xilD�������ϕ���5���4�1�O�Cr����7�D�����FQm�J������յ8�	E\ϳ��v�=��d����i|ܽy|84]��V�n��y���bRaء�%�]��v���؅�H�����/���Ι�v�1���U�>u!5$~�� ���|)�V���g��WU�]XXXRY�GQDm\��%�M#YBB*6vQM�?ԭ��&eY�t:r��[?�T`�m�ʣ�{��-�a�M��D����.n����������\n����bQ��]�v��k��Q���<L0�Ȟ����i��l�M}���zv��U����s�^,��0P�xgf�u�g�,�X^{(R���Ć�Tb#���X���t�������ΘP˳_u��CK#�mY�ln�eVZ��KAFk]�_������D�G�Q6��m�'##�"Q�Ѫv~�4	r�<�c���*���&H����jE��P8uF��ձ���iM�L\�@�������:~~A �:Wwy��QE��V����5�ͭ��Y���2�i�qL��l����,�_="vљ���o~[n�g}�qK�ٺ���7��w�k��yg/�Ƀ��ʞ�R���K1C�SH���a�H�C|ù�Fӏ�K��+
�rX�x�@�̵�a��󕢯ks����Eo��GM�7#�
���ee��O
�ww��� k2L��$�
��qC��B����f�v;3��1C<����($�v��39��?$��7	��f�Rq��'4=v���>�89�T>����#�7��S)��N����j��ӯ<E�Y�"�w��ձ"�K�����L�t�l9q@4�Z��L���^ͭ��l2���y�{���GL��殀�!�� ��f���.��Ç��gު�
�:Z;�v�äz�+@���&ŧ+%��ypFL8���_�gW�(ʱ����9��Ɔ�Ǔ��&�L"�/ʫ�6G¦��Y���$37�{�V��)G1��SD�N�GD���-� ]v��B�6�AA�y�1��-��H݄M#��C̮��W 5r+��-9�a��&�?�x��ChI3k�֖������B�H�?y[���d`r�v>�/�*	�l~���p�eh���\����}�/�#G�a�[[���WQ�Z�|ŧ6�X�M���������qѷ��ʣ����F�!w+��D�����.��%jm��;0d�wU[���C{Q0�������k��Y?o�4E�j���?#�#�
Ê.Wޱ��$Cc����x��{_���B�W~�5c�L�|TV�>��?���A���-cn�}(��H�&�����i|K=C0���	�<7�w�G����K��ն.�4�*!)7.hTB�ɬX@}Ysb�(;/��T���e����j����,v껑�x��;+�
e8��Q�>�v�~	1�mJ��hLX������br �E�d�nT.�:0�n��s�_.��@�(�#˨�L�,aZ����;G&��cmi<y�W±ygDǄ�,��ۨlI�8���y�G<<��7�c�V��T�G��j/p��u�0�b=I@\{���WM���f��`9���<�@K#�IjP�怸�2u(ax_��$_���,T������Ebߞs\�`'���*]8�1���$~�[NԷՅ�5a�"|SW�����{�Y��m���?�b%~ȋ���G����T��q�\���h���c̫��^�<ݎ_&y������Im��ӱrF� �����j�e��9g�D:my$�vy%�<�@�ڀW#�9X5YO�?�B��'��2l���� ����Bۼ'8��߳=��/rba!bB���w�Sܮ�Y���E�c�(��wRɗ �8R";Q�V����F����̛�������|�]�e�7�	�Ń^wP�DS3T!���O_�g)�<�ͯ�[ڔ�g��AKEK(�}2��m�ȷ�
ո�>����Ur�	s�"8)_�Ss�f7�i��!1��@ԑ��ꤵ{�9�[j�;�k�\��Z[I3�8���T(��2�BG� �Q�9��Z.g�[�~ F��*�p	A�^M�]�k#U�B1�gv-�p� 9)S�| #�D�Ǖ��R�.�s7�����_���������8nt������Xdڝ�ѸN�Y*T;e�{�_M��'7�lU��@��@m)
@z�!/"v8O"���@N3qw�
R0�'Uo�~��ISj�9�@�L��)��V}�i_q� ��&�BMc�dwb��J8u�}Q6�sx)��my�9)%%��� �2A��C���8t��X��pĂ�ǚ�����\�;�0���eD����e�ct!����ť[����"!�a�p����˾�ZUP���?�BG��P���/^�	^������ˎ�o���>�G���;y~���~oU�KC���+���	F�/��0O�t26�7�hD8�����w<H�lyu��g��aY[��C�߾zQ]�Dỹy
�n��>���,�]�$ լ�4�C!��u%幎�y�KtNs5~H׬X�'J�ln'�Xc/�������	LƳE��N�k?M3XXYIL.H*k�>�>8ұY��������KO��p��y{����Ǆ3���N��k�]�h*�H$�Y�S鞝�>��g?�}��0%��A"����1��ȍ����
G�P��\p�H��l���N���,@���mF8���*�㺭�%Iq�qX�fG>��bHJ�/���|k�E!"8�2�c��|N{{]W��Ϸ�ς{A�p�3��ո9�`���MLz�l����4-�~�����4��*�C�;�n��a���!��yɰF�!7(� �Q���lp�)*Q�%U�&������@G�'��Z�Ir����9��&o1��:V===�tx�`�6)h�������ks��R�DJ��lD���-n������I�"B�)��
	Gf�F����@�ϥ�0��e�E�c=�hQѯ���{|2������Z���|�t���SW��_gk«����cTN\�������[��fӴ�R�Ǉާˡ���t]��)v�},�Ő𮟃(?$~�@�e��)�tZ�)�##|�v���<��YOe8�θ����!�<<(�>OW��71�g�8��N("�e's�1�[}��+�O��ݪ���BH�+/��J�kktX�RRV&��I���?��6q8��/-�T�HiZ��X�?#�>Ր�Q������Ki�r�N�1m�p2��w�]aGW_e^�	R���������	��phA��+e�P�IT4���h�J1� �m��q��b��?���E����;����������ݎ�����ƥ}�_2�꽜�Ћ�TK]"���4�.�)j�R�v�Y}2�1�42�)'m��F�[�e��f�����y�~��fS���0�?��9���'?eS�޽�(&����*�<A����t��ݦ�c�j]�������M�ʍ0G�����#=̏����W���8B<eL}�����,���[�S�܀�G�tŒ�r)��@���G����ZZH�%_Ax޷�����<g,�|B����I�!;Gs�����K_����t�	qS�M�yc��dJ�6��'��_f���ד�������kn��eM=�p���O�tH��2�x(����v5���~�A��	��o� újcO�^�]}��fVWcm�/1=�O��"z����q��"���?��>n�a#	�T����1|a���M#�)H����Z|
�T�0�����~=��i���k�8;d�q�:=��|�eM��C�ťd@6��l;�5V���Y��&BB %�S���f̴�'U�ub;�]�p��o���<���t��2q��2��y$�GL�=��7wo��,���� R;G=���wZ�夓Ux��R�C�]Gj{e[c����� \IS���|�4��Hu���tn� �7�4�y6)8��,�gf�&s����N�Ly%��qk�˃o�뫝�{@A� ��Ae ��ys{	(�?����;�{���!���@�C|q�c�߶8C<��S�[Fzn��Dw�zR�f!����U��r4�Z��m�jªk�-F��j�k9M�h�si�q��.d�$[c�q��~��M�u��ưcl+��A$�xtg�7���H� �H{���7�?;�ipJ Y�J��ݵ���G)�u��%-�^�}�Ě֙�`�Ak^o��)���d4ٝ������״���&�Q�'�sT�9D��������������g+++���X%M{�c�����7]߶���t����@/V���$^��n�ԑP�B�ԑ#� �>N�Y���p	AR� D��[�[��O�.�ݝ쎿m��%�er�bl_
A�`��Fxn2�ͫ8��J<&��ql+�ް9�ngLS4r5�K[�H�9�}�i�&�.���k���,&D�?#p�i?�R��#���Ve�}���"~$_��R�0����G��B���j�\�J��O�K��g�:&�&c)�Y�u����\F�#^uZ~J�{^�������)���م�a��d�C7�r��i'HO�&�yb�CP�|��.U�� -R^Ja�ՙ��6h�����K+���+*���ϧ��j����W�!�O���}�Ƶ� xrt+NW���}�t����+�W�%H���N�ir8�5���|��?�ND��35"hʱ�>Lg���W�ꔫ�5�,&k1n�B�޾r��\ě�ŀ�v�u�g
�����WRc�O���f�l{P��d
۟o�^B�Y{�u�a�r:���)�����>����x2�pz�q��)cy:��8�,n�0�T�5�����~v6��:��O9>�܉ѐ�[������$�/7�����k#&�H;"��	��?��$ٕ��8�\���?��� ��HV�k�Я�ڽ�~>�zi�yʻ�qQk$�)��׆��P���R�������-tDv.�����KB�;)���C�o����jx��	k�����`��������� �ϟ%�g%�g��[p5�Q̉���2⢚�� ��K1�����\	.^��SN��ԩ��]��iI8>7���`��E��� �4�ӆ����~i:Z11j�����>���Ժ��8'fS�U�p����T�)I�4���>z�Z��M��W�a-�Wc3nt�ӡJV�4����{	���O�b��|��txx���5�8}���'YY�_��rX^�!��tx=kN�5T?I�K"���� ��]Y�<�76I��~��R9
��+���=$y/�Q#�Z��_�ђj��nU��H9t��E�L��r|`Ӹ���ȯ��A��hUARŶl`?��,��K�s@PE��?ˠ�평,K]:::i�uM<���Kؓ��`�D�q+\���=�.�*�M������IG�P�e�;l5�:HT611�X����`����b����*�(�e���i,\z�DûStӼtv?�[7���\
ޤ߷��'`�_(�;h�N�@w7��v�2[��H�r.� #T��=��_�Gi7:砫xDh�V8�do~B�J�٤ّ������c�W\u��12̯�^�0ҼZ���6ӡ79J�j��������Aˑ\9���|=�^e���-��?�E��fw��-�j�[К$�=��������O��r1s*	�A��@������E��pO�Z[O�Q��lʧ�$!��z�Q��N��n{:q�JA��t��4�hV���XTS�6i7���E� .zh�;'
�V��rA��P@6�����' ����o����B��H4Cf�;o���vOkn�Δd�����F!n�� ���#��_����h|���|ZVt���TI��k5��`����|Qġz�i��E*�Oă��TBSX-�,neA�ջ;ut�Ὣp�4m&��)O$���ON�o[N����IiB�LH��k�"�h������B(���ۉu%�BEQ�y�>[r�QNS��>H�V�ѐҞu�֔I���ݷ�BC�3�����@G�J��q��]�hѢ$+�K�z����eܛ��a�@�KC����{6�63�2��{���cI�|%��Ve�lF�7.�
�(i��MF�s�s���U=�e�����/Up����l1�����w]Ox�^�[�fI�p����_��%M��ŉ��|�*�Բ���v���ޓ�t+2KӢYY����]��X2fͅ�-Ț
�琿��EpB�Ϗ8�^��ʁ8Ϟ�OL,��u��������qWl�\)�cs�D����v��T`*���B5��ڄ��`�����s�M�Iȋ��:O<������a�)�t9�hQ�Q�x���U���^RV|�ld��.�d�m'.Os�}!m��i%�o�GK�����k��Yz��{���LH�=�@bb"�{�N�%�����_W�u�jW�P��X��o�;u:�D�T����GP[Nl�G���.36t��L��}�tPiz�0=����h�l��X1���`ݞ~v+%�~��u����k��r�6*:��=7k397��g��#�t�A���^�� ��^6~�kٻ<���(f����8�?�`X�0w~�G��*���H}�?hm�Ѝ9����i��G�R�Y�|����8�1��+t_5�~oL՗>��`,;�m���p�lϨ��?0P��2v�B�X��6:t?]��KIS!Є�_��{i{��i��t3�x�#d&@g"@' &�[sʭ��ҫ$�¦�����T)E~�ٜ���'t�?�\
��qpA)*F�֐����b��lp�T���j�o*������V��_��5���Sd/�]j���;� NA>���-
�}"�I9�w���]mi�\�3%�:��Ou"�X��(���n�D�a���JZfA-�0����~�F_U�1#�#���҇����u�J�m��A��T8ƪ��/��@x�|נ���遵��d��Zdux�G���U}�2�*w�δ�$Z�yZ;%~���؏vL�{���7�[�:��<��H�
�j���Lc����kge� M�����vJ����r�N+������+��F����ⴻ9]�.�Q���QM[s��Wu��7������~�g/MP�����m�y}�l�I{FH��N�0��a��
�`��6v�����B_F��A�<y����Z莟��-�(�RjgN*��'��zhQ�[���A1�l��=���xO��;\k~�S�����}X��ʍ��Mc��F��y����Vҏ�����=`�-=?:��5u�;N-�G�S�5���<
pu9n��o�HQ�ǰ}|�ԑlbb� sko$�p�>?Թ���ђ�[��æN�������k���G��y��5R�8��_�w���j����+Qď>�վ>D�牴M'Cbo�_��I8O5ܲ�<�z�yO�=+���`F�����!ANz1�h�2����S������8$г� -��V��.uO�Scz2�46b�a}kO�1 (l�;� м��{�}�;	�2F���X�t�ccA�`�����s~f��?�a���я��]�Mz_�U�A�k��݃��Cy�2R��3�>�^`�`s@x��p���ۡ y�h�u{�*h��<����4��kZ��<��m�lX��8��/�:|�@to�N2_X�S?"l��tZ���y��l��A7%Z��4���iej�5 �l���ȼ{�#�p-�褶�(F��;A��I��<j�!�$	�8���^M������1Bf�������QE'��1%�5�=
V������:0�P����s�����������H?�v��fHԝv�F��gN�;�F24du�ɯ������&�����*��@⺟ݩ�J3� l2�Hق7#�۟����1��	���_
,ZK+��r��U�O٢P I9�[3���"�{:r�dzd$�z�-�im�a�f��G��(RFNFܪpM�j"�����J�-rs�}K�[>�g��un��еAc�i�鮷����#� e��]�I���#ȑ(EqJ2�H0���؉.Dc{�<~��v�."n+?�t'�;�\�ID _)�,�A>D����Uʃ=y��E�q{�gqZ�o���qA���b���'�w�^N}�w���M����Z���mf��Y���{�\��Hj�x��3>�U?��pDGڕ���t,�s�R,���Ql����=�h�O�����O�b�Ë�����O����~<�D+>��Gx7r"B��^;��l���;?Øy?j��>�������Ł?�#>�v��*��՜ ���^{m��t��C1�n�G��jUdz���Q?�#3X�o:�憮{@��ų��[��'=�j�P ��F!��ɆM�-�Նg=����V��]�5���"�i��"�zh�㰷�PD�U��Y��3(P�� 5Ŵ�={�ޏ��s�.g@�Cq�S��?�Ж��;����}��hJ�jڨ�r�l�����yu�|ݧ�%��k2�0�u�e}�f�R}� ���O��_�.@�9^�=�b[�ojv_t�S/T{��Hh>�{�#K�x=t5f({��_
t��`���u��Ħ����7�&� 4�ࢉX8!��;
_���[�,������ܲJ�W�y�)S��.�G*cK�*�O?v��f�?�-���F�#��WF����+e�-T�
�x���7�{��Qn��_���!^OӇ�S��S�3��AJ��ښ�1�e�g�3����9T"N���xl/|��v����Z�8�>��������g�{�[�fE������?�߄p�� �U��>�JY��2�裔;��[�vB`jNb���M��N�a@D/�+QI�l�_/Ev= �8�a�D[��v��8�����(�{�^�s����>��L�=���Bx�%�s�"2������X��k���|������i�������Q2l�_u��60W�3��xR��Z�R����W�G���K+bN����;C�jܖ��N��cy~�u`5~_�:h���ĆH=���Л��x�e���U*Ys���A�Ʋb�[���ϛwYz�~�������ߏ�t��hgp���F֗�J*Gb���J7%������������� BѢ�����*sbN�t���b��*�;9Z�ܸ����(�+.C"���LTR�>/��k���L�/�J�ĥ��3���/��-k>J�$~�d�Y�^09��������X�/��١Ό�l(���B~���9���m��C1��#�ќ�rA�H�Fp.%]�s3'���vق�1�������J6n��~{�*�)gK�&|a�u���㗔"�$�B�d�z�����>}����������<��� �R7��iMW"Z*�cL�t��Щ:�IK;p@�0��Z��)_��ۓ���az=�Ee!@;JI��K6	7r����Y�h_F�������NJq����i@���,�b������Gٔe�ЅH� |� %b��E/����.����4ػ��|�'d��q�ܕ��-ٿ�O��&�&"�Qb]{`��h)�����.�(���Qѭ��5dF=cG=d��A��i/���?�c>��=v�3ߊ������Aj���V��<t��ʖd�Y0x�?�S+��M�};I�;L�[�)��|�?W$pQ��خ�+��_��E]��w��9�.b8�2B�A}�u6	�A�?6�&�|`�/@N�EO�h �o���GF��h���:y�W�T�H�Sض�;<��X~u��cV�ȍ��	�c��|k���y܊�"J3$�%\��C2��>-�eL�eQ�`�CD��>q��[�x`�7ʶp5�jD$m# �'EQ������JqC�`[�~�˨P6[�|��b�F��B�l����_�]�
�O��N[�BJ�g��Dl������IgΪt�a����=��v�wtAz�DB&<�*;�6���(�U����]�t�}c������Vj�v��#��4�7G�bC=]G�zKt�������г@4����o��;��	���� ���-x<!ҥUB��%��� ����:���BuxB�JA��4�qIϼ֑���#^�����ˊ�8^���v�Qr,8���K쌹��zOu) �#3R����^z��G��g1u�,�>������~a�Nk��mO��z��UW��E.�ГN�i�'xm��<�K�8�3=����k_4���d^��mIv�����Fk�{���
�LD��cD��q�3����`t{��qwl����[���M�Wlt�3�6u`Ӥ��%�o�d��� ��D�7���qZ����kGk
��V�����~x��r`R��ޯ���'��|�g9oP��׽H=mn@�M�k�ǯ[kV����)3����̍e��q�yab=(~\np_L�|)��
����/�S���<�l�:��;M�x��$24�9d5;ӱ��=鸊lB��vsY��ieI8ׯ�)d�֔	�L�ڢֿ�؈�n�A��%
���T�]�G�"lK�D7}X��F��m�ݼ^�IRZ�ԘH��4�_i ��珤����>���cmտߚ'�[7���{��[˯�lY�3��F�Kg��؛��4x5i�rB�q�/[��@�_呡]�_&�^v2�ei� /�<(+	շ�4���)�z���ٵ���Y=��Q��F߀�*	���.�l�¨��D�����O=����5�@��9Lqp_&!���[����b��%�o�n�e�	@�>Aw��w�#^��,ʇ� �i��XQ��l��e������b��pfp?��1�6�v�C�v8�����H�*�oOK&+����]�������`�R9�P��]���^����F	L�P�Aז�3��$ �"o��#뒩��n��u�������z�eQ��r_G�v{��	��g��)K�k�x��g�ܴȳon�c������6��]�n�R�B��S�ȔY�d�k��ݑO**���G����#*��2�cW��R�2|�����U�_� �بwj��4�h���9)W�"*46<4b|���j�j���O��ȃJ ��Cդћ�p�5ȍ���=������y�lGf/U�~�3�9��
����%���>�r��iT�?�u��IZ�C5�\RN<����	�_��F�e�NN1���?ၭ�Y�հ�;uv&�S���E�(����Ku�/Gӊ��zK���{ ���Nd���.TA[Q��R����.V�獑}��!�G�HZ��a[�&)�������J�twit-B�UF��v"%����w�<���&��T��H h�Qb!��
�h����k1à�Nh��l����q�s���Q��Au5]��������ww8����<ww�����������V�(
6�g�Zݽ��l��gqN]>��E珡"��9}�2�Oɺ�$��F���	��&X��Kaq��䍈Ľ�ŰbR��~����)���w�'����1�KXs9�K_b���8]��9M����c>��0Ek��w�yt��b]���W���aq�R�Z*�:��,��H��u����7�.����t����?���A(W�R~c\��h��0d���_z�s�CP�hEgÈ����o�d�mC�mE�:HYǁ�����]�)�"� BE�y���lެ��񎛷U5�iE½�ݗcힾ�&���`�o�+����LS-� ��G��P�yK��ܼ�A1��H�9�oj���0V�{��� ��e�u�xp�����6g���W�ߧ'u�p�NOJ����8��n{ܸ{&��r.�mق��k�l�Q�X��ꋳ���<m&@M�`1ĕh5�!��:����FܶfZ��4&���_<���U��ID��x����V��Lɋ�S�)ّp׹�{�lj���`[���!����y���#x�O��}/E����3�1�hMAǏ����`a�{w�>~2�����N�zz�9h���7��
�9{�8�Ȩ�u��p�.[��:x]=f��a��8�� ���*��W!�Q�x�R�������"�f(eF�U�(j{n��B)�^J��//��$y�I�N����%�'n߶�X��
/��&����ܮn�z��w�;*M507L��X�՘=�W��K�R}�\��GOTy=�����B
%\í��Tl�D���v�-�H�T�'�:y��h�K��K!c-�=��aؖbT��3���sYW���O/�҂��>��!��2g{���(D��!3!�S�J`��)�Z>SCy���of���N�����0&ӡ�q��px�!��袜�=�
�n^L�-�׮�Y��>2A��h����Z��Ԩ �N��Gn�'zp�A�G�
�CO�Ύ��d?3���}OWt-`�~�ȕ��;�SP�='�c$&"�YSґY��u�����$���S_j��:?u|�$�'���{�Q#{�{{DP�aag}�p�O�f� V�����#l��an%8��X_ܟ�p�J��rȒ"#4��<�m���`�F�D)�Ŝjw�S`�D+Pg�_T˨R�h��T����i�K%W$�kZ
+�+m��QCo�S5}�&��33>= z� �˘b���{��	��;�q���B�8R&W���D��JH$=�p1����֙��?����s����&ͼu]dW�F���U&NNum��n��Hx��}R��T��ߦp�f��"�@��.�J��uh�r�j�b2������E�kA�+�šS��bR�"�Ӑ�H��9��R%��6��Yb��9���E)*e��眜++/���X��mr�g��v�"��$���[�C(�?�
�m������pZ��dz)��ہ9����P�FQ�(Ƞ�)�=-�/�j�^<v��D��0[C>t!��;��vnn=j;��]�l#k!E"F>��8�Yl��G_d@0�GJ`�A�6`a����VO�w\o:-ݑ)�ȇ��0���]�υ=�Ή$FJZ����Z�t���������0��S5О��)�ٖ�!���x��;�g�|%�׍<X����Q7+T7�O�(��;̈́�I/bX����G�8L�pDip��<0�^��HiC�a2^B�H7�<�L�����~�6]a�=���h/�}�xq`�9� -�Wި��9��X�.t-��|$�1��n^� �x�<��()��ڄ���H/0k��.;��G��eq��i��Zq��$Mr��3��xO&9ݼ�,��׋������ڜ�M�f�Q7g= �9K��i�Y� �9���H�V���{��O\M�ev�]O(tP��-r\l�<E���k��#���Y�����n7�jj߲�,+���^�k!���'eG���X�A��bR=Eu�@#O��;�0*��W��;}3����J�`$p���y��r^�)���(�I?��x�{�o�{�&`Պw"̓͜��=���'%)(�2?b"o����'���cCK�o��#o���v���+�k-J�Ѿ��2�@5�)��-b�ʑ��k`1��ςRCEF6҉^uH������"FO �M"�����^_��J�<���� ���'��t��hҙ]���Bg#�Δ�یa;��0�=l��0O���Q��Ӎ��QF��GI�zC����K1U��z�����kd���C=q��RT�ftm�׮3���0iY7iX�qi���Y�J�"z쟉�o@�_��k�{|r<0]�������|�O���aN���5�{��{�S����ӌ+J@�Ŀ�&��Ӄ[	+U�ʤ�l;̂�%�i���yW<<��vf��fd��4�|Y1z��$Rk1�uPR+�,sLEHz��վ~k�N8'��K$����L'��z<��p��0@-�b���}�i�fĈ�'�1Ff'@Ԅ�Ժ|K�d���TOcY�T?�{r��~���ЭQG���Q������/�y�q�h	�`�Pm�����J��7M�
dŞK�J3c�2C���ݽ��i�u���ݯSGJe�Tf��a���GD�&�g�u�h{E2�#޸��k���p7���AH�~$e��z�V�H�����r-�Θ�5�	B���u���D�C�Z �� ��LV��>�I*� �E��^��O7/��~eDV#��WhPLHʊn`k��<d�	*!��'���}C�v�X�f��(R�;H������e63w=�2����0�Ko�h~�*ܡ�ڇg�X��EMi�/*��6�TZ��c�&�,�c�*4*t�8�>Rqx�wwn4�r������^t����VJ~ۧ�=C��zz��zz˧�ss!��E��X���,8������G�#�P|C��da���
d���$�a`�8V���A�H�> >����eۦ���{�����߾���9��zpP�Fb�,��=����
�c��`!�{0Ib�o���y�`�C�O������[�>�\��RU��G��Q���b=<�-�[ ���CE�9��*3�r��x��u�w� ���&}���4�`�\޳�
j�d\SDr���t��U{�/,�4�8(��xIgg֛�ۤ�4�4������p�ܩ���D����a�[� �&U�������N����ۦZ]h!T�#!�]�f�s�@��f*ÄM���-��:��C�a�����qS�RT>ڭ͊���ح���K���`���-���
FpyEELf�����:��8�B.��pl00'&n�2��D> �-�ZIBVv��R`ai����m�۟�������߀QS�'QA��0	��+�I�f7�?���]��jlj-P�蚄h��f�2qH%��i����J+%�_��h��ҒT��w-�n���E���v�2X@����Ɣ�}�F���cc�-,vc٧D,,(=.��&��������+��}q��V�
Á�)�%\N=�����.�l�1(��h�$���e��{zi�r�c��[���T����8P���6hX�A��h�B�3z�OB��p0���ƒ)W��b����8��}�#�Ke��dh���S���E�.M���;��̨Nb����{�U�Rȇa5T	�Ϙcފ#��-�e|�tS|����>��Oı��b��B���SCi�z���l����X	����4s&<��r���/�A�,�؊ߚ{wA�ȗ�HZ������5g2���䈴�	�d�,��������g�5�J����q&��UP�"�	.9i��󒎕��F�v�g��47wdg��ܣ���p @<e�9�/["U�|��Q+�ӏ�fH�_ZҴ���;o �`��n.	�ʙq%��V���� �΀)g�3��x[X���>�%��~V�C���&����>�CL�`v���?o$\�IbRR��?rY���/�>�M�*C�!�o��=���&x��b�c-�ۀN���? ����4�/Z�&Z��蔫Ľ�K��ǭ����4!��T>�e���Z�Y�iW�:�r<��x���|D5�0��:�,H�ϳ�$�&ʯu��`���w�-Qw+����zQ�.FA�>!,�\��s����i�����?t�5uJF!6阜�$z�a���>�뻌Q�NL�*D����*q���r8��v����#�Q0�S	����� ����0���U+I�/t�������0��{�zЇF�)@����8�Ͻ�:��s�i��2fT>�Urz��T�	�?x1N�i�P���C�p!���n2]������Ep��w�����r���Z����w�Mw�'� ��X���g�zs؛��+��M/��D��x!oZa��*���⧹��E�~�2k�	%��eC�#��g�Sݿn�؆�r�m�͒��>�ZH�y��LV�3�E�_H����K���#D�4#;C�@b���	n���%c ���1k��G��WǡC����-S*J"$"�ʫ�Dkq�!!`�oO�S�k-'�< �ɡ3��+}���JdXN?�˰(v&b �_%��:��/_�Cӻ��*k==����/��f�#���#|Qȿ-^���O3�0���) Bf�&�����铼vJr2	Z�Ԉ���}R�� V��&9�����G%w��j5_�H�L�G  �.�}Z݁Ľ�r�A���Dq[@��b��MV�ͯ��$����I;9�jzz��}����f\ap~9~�&�(�!��x߰e��g�vn8��aJL��Pe��AAl�)��H0���x�6E�4�n� �������n�N�Ċ!��q�5��x���瘦&jVV4�د5������x]�nx��(+#�d{�mb+��i��Bv��t��Q�u��B�ai������WՉ坻ǡ���=Qm.���e"��L�r��i�
 "�U/�iUi;���>��ҹ[�/y�#�*Z�
S<q����6bK�na��A"�{g�	����{Rt��G��R���	3���<�<�a��_w�?���+���9�s�o���O�cf(�ĕ�Ϳz�	 ������6�#�N������d��������ԙ�:`#�[ �í1 �TU.jꉯ��Ӏ ��U�����=3c������6��=��x�W���کc���$�}�9�����	��d�6rp�>'�{�D��K
M�u �����\'3�(��@�Ɗ�"������*jh � �J��V��-{�U}��	�~�
J(AQ�����E;��0:؃��/�j��&�=?$�d|���` Ȋm�»��`X�.%�
<4��XW��9��Z��@� ��/��׋I`5S@**	Uz�u�S�����=:u���`�`u��dS����X��<nG(��lQ�@�$]C]�[1�>��H�ZMD�/��s��ԑ1�Wg��B��L�@��o�ݠw���ϳSsIܟ9��z�=5	C�t�6���H@��v��q�aՈ��x�l����f&~�loE	l/F����m+"�p���HB�~�/�h�h��y9%�Je� ��əc7k��o��~���#Е���oW�1����۩���o1�����w��F��r��^�1$��x����fө���AHK����i���ɞ��V#|����W���m��1<~ӵ���#�*�4,!�pZm�LO?p�?������ɢ��/z٧BONN�7�̼)�c��,]���=�	KR^��S��7{���ƻj��&�e$y贈����ۻ��ݷ����'�z���}� Eǩ6{h�!p�s�}�`1�"c�f�IHS��k
/Ԫ9>�&���q=_�
�x�k_����� @�X���h���`/�`�:37��:�T��l7��^�,����)qab����zxx������Q�э����O ���)/瞧?��|p�L׉�ҌFR
��҈
2)�!؈�=��$&EY�Xs��m�khh��d �Q}CC������Qeઽ�"�,�M
"��6u�g��V� �?r�����p��Y}����N��w/�}��������"��5@��蹖����� .l�XlMC�;�r�a5q���A�S����G2bH�<���$Nʪ�{��ɠ���.�%a��n��-q =��A�wn�H�O�VJ���,�ͭ7B����8(��s�g�Ň\ǭU�~?8��&�s�������wz����Am'�ݕ�A�*���&9�����-AQ�={IW��F�x��S�����+��a;�Jt�Ӛ����f��i*́�8�	ŗ�LQ��y��}777��y�=6�L��|�S� �g�\/�t<���l?�Kg�dt�eIJlRi���s`��u[T)y��j<��PWд|������
X����Jкc��ӈ���>��6�f:��Q����;O�TwŲ�N���s�[~��-���ϗ�p#{W��l�|'���!��(�n�_k�GT�ȠF�
!S'9f��i���F�	����xJ�����ޡ���p���h���W0s�֓g�G�bj�I����5O�>ٯ�ӓ#@�g���/�z�D�o��p���=��lu���/�>�1����.�� 2��zT�&d��r�i��?�X
p��{�(&4�U�}���@��I�V{�~ݕ�IK&W��M�i���z����S�V�ˢ ���C����"N�&Z6�-��!�zeT6_P;�P8��+e_s)������y"��v����ڛQ�A/2�}�a]lTdA�2t�&R,2����@���`��9����:�Yr,
l��-��i�`�Io��^ހ�9�ج�`^�E(����\�����yз�,P���9?]��m�� ��)�qo}M7
��tDT�] ���#�����y��8~/��h=�m=m��U��~|���g�E(�X<.��7�(6����ρi��QZ	��&J��Ȅ*�����ݏ��f]a��Uf"��o�hã������^(e5L)��`M�'&#�G}` ��z��H�jKO��@cc�9��
��i���ݸ�'�(�x��������f����Pl��<����m�������͐���f���$2ז6���|��w_�������)���.b�ˬ���S�u&?"�^��d[��{��п&&4|-`#�C��Pe�t�A�1F�����F�|̳�{�����)-��+�����>� ���`���/|A�^���Q�"x����+�/]u���YaS�����;����L�tb>��O�Ӊp���B�����ԟ�I��� >��HME�W�K�8�}�U�ӋI~�9���,�m6&@V�1��y��=�'�q[wSM;�)�ª���k@QWP	��S���}��S�X������3�F�G�SMߟ0b��vE��bD�̞�=w��w���	5+��@��x(6R�ҽ�ђ����G����39��|{��c��W�8�]2�z4�V3��b1���b�&r����d�����jNk��އ.MA��D4�H�~��c�����I�+�e�.�������y?�8VF�Ī�]��km~H�F�Y4��e�._��悭�h�o���csUU�J��z�l�S>�_-���χ����}"BG?od[7�.4Ұ��?6�r$WͿ���������7�9�+ʣ�����؅��h%%%�N�n|&��z�ғw�y\��Pk�6j�,ԛv������"�h�g�j� �xq+_��܅G�*6���
�o�7�|���&�4kj�ցl��}�@�譶��㹦���1��%W�~�����X�ןy���D�u���9�h��W���V|��Kn�$X�^匿C��\&���b�2D-����%����)+�x��㢔>�t#��L�ʐ,��5A��水�<��řIz�`_�XuI��%k�?�>,����z�}}
	����<��K� +����l񍝂B���N�t��3�	�: ���zM~@ռN�Z��G$�߇�
�{�o\�P��g_���f�"�4?O]�2")�{�B\e�9�Ͼ�������@�D�������G��c����Ra9�˪*-ڗ� P[�r�����8�A0, �컦BG�������V`\m4r@�6�o��m����,"��A���Q�t�x����甎lT��zI$�N�:c?阻}@ �p<���n���Ӳ.�����2����C�[U���֨�j��z�������nW�P5��`�	���!�A��k����!_�{��Y����R��������ŋ�/E$���/'����G�f���Bcf�%|}}%0�>�*� M^��$��Z�,�Q�R^��~��;z� �sH9�mO"�l$���3@Ì�SW�j$"���|�I�A(A�%my�<)�bQ�XR���Mz�⎇��ǴK�Rpo��k� ۚ�2=����)�ڱĔ�\�]�f�W�@��mn7=j�B/��[��"����C�̢������"���{�?�4@>v�2�Q�^�s\�l��.��6	����ύ{|�nq}��D�ۂ��Z�qN�}�&�B��`<�Pbo*9{]��激~���~���/� e2ʈ�<�a���{3ذw}�=�Õӳ��SBZ�Ò̌�I��*��U��d�I��(����*��en����\|��]��}�B��h ��4*.x�:&P\ٓv��)6ֺ��MM}��47�iL��5�I�0/�(P��(�y�j��3[�+K&;�	y��Q�Y�f��s���e9�����An��N�J�������y�cD(�ň����%4H#���\�rc�O���6�pb��!dY��34��6�;�ï n׶��#p���QL��YvH"�k ��b�Uel�E+P�00�� <y䚿�v ꩗q���7���w���ۮk�D�3$�0�Fʬ���.�g&��$s�0�����ŋbL�D8�����`�Fx�K.B�㦐DMgʙ �,���,,����T8��,�����bl����|P<���`S�����ѻJqqqTʌA���J�����OebA/��v�h������߾�1fO�Ǽ A�T/�?�u~&N��&&�ڊ�o������y�����if������h/��&�s�*���9�g�nj���Q��V���i(s�뺈��G�����#t�,�2#u*}S�!�T��**��jk�E�ἺLP*��o�
�'��m�Q��	ĄT=��6�iT���v@M��Ľ��$����w������q��������,?���v�D���9���j���H
��m�m��z�n�����q5�����NN� m�Cfz�/�歯ӭՖwb���f�j��:q3O@�JrI�6/�!c��;b��L�`� U���q/;��8�h��IQ� �k�P��{�-��3�پ)��a�$�]w"t�LP��d#�W�ѿ#c3�E�'ĽG����zq����!ٓ��5v�����פ�Kaһ����� ���?p\��������쇃}�F!�.�o������5qYڏ����dIq�^I��y�������6\9��� ��X=�M|@lC���Ho�-;�Q���4:������.o������L1����b�y�#�:Pҧ�ab�_�(P���+ʻ�$S��ka����U=ڭ�ɺ֡�a� �e�R���M��΢LE�1��:��%����Ye��,"Ft�x��G6��1[H�U�#\R�Ae���zø���8���7��g̨T�K���esc	2T��#2��u@��ЩK����� ��?c�@%���0w5���_��37�W��<q�m�<q���\�j|Z�EPy>�K!FTm��w̿��2�&����U}����~zV���q63j�ngLF4����>(P�q�m��B��5U���h��}��w��7��i#�	i$��gڻ�<.#F�t�j��oGsXX�D�V_�|����*)[[:
���1!�@�\ArL F��l�h6E��C<=�§i���#�u�ȹ?�O��"dq�|O��!�]p��S����i��'ٹ��˯�B�:y{Q���D�ԭ�^����p²��@{�Ah��o�9� ��2!���%���W`�Ly�h���)��և
�y���sUk=0��yy��v�wY��4~���+�>W�^�`�Q�퇥�g���|�������k�;�����G��)����m�w����f��apG���[G�σ��:�J78���;q��B-Bh��b���@���K�@�Q)0�Ǩ ���Or�]��`�G��7e��
U���������_�
f��kV$}�A�U��R�O�u����e�ތ������Σ%!ߩ}yub��,�3���X3�����,���M���`��2����i�?��v��Ng�����3E4AM�xn�,�lLqv��D�r	�cd����g����~x��ߩ��"d��J�!�_s�Ч��0�C?7V�ͥ�}�|�}-�M�Gwx�į������G<c�� ���ϕA�	u�Γ�D��ǀ��˱�AӅ4�eJj&�[+OLΝ�aL1�Q�Bp�h�	���5fG(�������.�i1�[� d�����IG­�:jnݮ"\����j���*��v��Z���Vs��u���h	��Xq�06�YX����P%�rxG%��}nƁ7�y�0@BKkۄ$����ƫ3��ο�,�}�7�9c�1�h���������H��I�Ʀ�-��Ն��\BvI�.\F%{ޕ�m�/&@+&�[����Ä�����3�S���4ԚG�'�H�J�Y*z{Jᶑe�C�yˬ�?���aB�#���(P 5��:�Z�����;���S�o���w��'	�B�g�V/>�jx&�r;��s��}mӧ!%�F�����_��2�I)�,O!�Ø�S���
�m��m�Y!�Q�������#f1a��бVx��sݏ7�whgG9)�}�"����k��@�^߅��$#��fa�i�G�*5��>,5b���- �/�Z��� Bd�[2/��Յt:6�G��u�����!6��)����a����ȹ=.r�7Ң�r��R܏AW�Vl�v���x}��V�<X ����=oj=���5�P���f���}x���5�	��~�0f��BGg�gCkҍ�����cV��x�Y�NM&��D,+ns������
���������2��:��j}�#2u�D�p!�c���|h1���L(�}oz�pA��_�����T�o�c�+1�+?�6T��Z���;i������=p����'z���I�0�LŇ�(��n�Ѭ��D~�B8��}���;����pE-�cW�uC��c_�L��J�d���ggq�5������*��C��XX����<�mJhL9vk	�����9�&(����J,
�����A�_�����{��6�b�OL�K�v��>��p(]UB�8��=@�}k=�[ceQ��=� ޙ��l��V�ˬ��D�Y�����e��=+����1�Yz��~�I�W�p�RT&����ȍ�
��,a���`Y��@���*�id-D\��Bb�WH���=@��"��e��A�F⚀߃y�[�o�_t��pr��VV�~Oj���$�Im#^�Kw=�8!��#f[.C��ʾ�������.t��-��E�>_���c,�G3I9��N07\�a/��}5R���E��a6��w9_1�;i�m�?=I�q�u̸1�xo{!� ���Y�ppp(\U�>��dg��|��Z>�5~��s�i��د���k+�x���������'c�p+)�_��s}���:ͻ���uhli��&��Ug�>]�/!쑃ӣ��~g�G�#�������Bt1�4`���?0��:������v}�Գ=�����f��C�v;�X�@����Eb�3��.���U�&N���+����7frc5{��`.� )�~'�ە�&���By���W3ƞ��ʝ�Qޛ�S1J���82#W�'}IIH$����ƓY��P��`��p��ק�Yד�
����v�+<�j+����]�Q�S�<+u�a/:�XFj[�b%�aJ3�kO���SQp�n�rn��W�H�p��c�B��䱿�ܷZF�8W,fi��W,�[6��|��,lj�<W�lY���S�>)�p��B j�{�	i����,v��z�y�q�覆����b�i���@/܀q~D�������y�����֤B�K��ߩB�y�,L��^��[�	��|�OJ���K��B|Г9��H�%�4�p)��f�`Q�,�HW��#�C�K^Λ�e�7��'gtV����_��I!��c���?���a�iWi� �V~�"E��u,���������q�z񹫯a�(y����~��n!����d�ꨓ�������2E!���w�L�
���^1E�\g�0��ˏT�	�`�=��Ǌh���[�S=4�S��J�t��tDS��4Oc �NnH��u`�\SɜT�V�X^�F�z~K�n���L�`�qp��V�Xs�Uv�1���$�K�r��/�R��RZ_qUw�.My�Ȣ�Wq�?\^�YU�*O޻��;	xs����,�oM�f�G���8]1آ�����)���}�^
�о�G����T��qr]�{G�}!OK_����Z�O?/M��PP�c��^g$h{��D%F�ϗ�@���Q����khh�LR��q"Q�˗8T���;C�c�TZ��6��{9*�D�}��� �M3���Z4��lG�������|2ߍi}��}F=�=��T�(���	���4����l��*�W˕k��w��l˻���2����ۛ�3������_2\����ڽ]���Gv��h���O�`1|��f����AA�A�ʺ�eB�$�ŵ�^ ��}s-���(��:�2G��Ȋ�7^����t���S�qbg�\
u�6p��_'�e��塿?�UP�z|�52��+(,��� &Fy�x�f|^^^�}�6s�ɨ>�8,�e,<�P�P�S��ۉ�����-PO�L���YO4���x`Udw�=��JQ (R���Cs�.6ڀ�R���}������u4m���S~�ލ e2�Ď�S6�j2`�	�����M!��2h�0R/t����7[!����_
yU��i�lMu���x�j�%Ca���&��o%�xuֳd��.����i=�ξҼ|�)y�!W����K�CG���EˍeJ�?�]�6"7�/v�3 R,��&]�&�"������h]��~�z7!����`M��I&v����-����M�^b�Y�������'ߎK��u�q�I�I��r�IoJ�9p	�_�	 7\i�̯^a'��\dk���g;
R��f���|����H��v�ʘ����óxȹR��՟%U��K�㡬�@��+��#�����c{����F���������F�K%T2E����V�M%,��ԅ�_�'��f�h�ZAG��<�al#�Q�/m~a�C*���$`�ɾzp�Y;x���p���C`:9���7N�_%�I��a�L�"1�Yp�Α ���X-d�ʴ&։����c��b�;���>�.<'�\�"��J�Yj��	N�Z� _�%6�_���Ʌ�5���!�Yij��h�L�/�nY�͜N��_���i�D�X��֦�0+��G�\�z�N]�N?������󉳭��sA�fr�R���>��)���Mjf�%�?�̛i\K��y�AO�Z;8(v�
�p�
�����9���>�SB�l�~l΀�45:D><<4V;���@n�v�M���7�P�����䃖��]�ۂ��_0g�M�n�7������ݹ[�,��D�z�Z<1�Cr�s����bg�Ŀ.���`d��$"�R≽��1�,�cN�t'�HGb��R�^��(���󭩘J��#Ҁ�>]-O�;ERI'���L�(��&���CK��z�G��ɟ���'�M޹}~fVV`R� ��k]�X�*m+��jy^O�,�N�!7�{e��	�v��؈o�I�w��`^]� �Ќ.��ʴ���d�z��z�a����*�Nn�Z��Twe����i�����s�vQ�hȒݝ�F�`s�;;}�QV��EI��B��y9�u��s�P���I��������充~�A.F�4���CX�!S�8-g�Q���8�Jԣ[/��IW�(�J�Q �vUCϭ*��$���ʐҷ��w3
O͐1-YWHǏ,�	�0P�څ�0���b9,�x-N�'ЮP��8g���̲�zuy��+(���qn��w��^^��ZT����O����)�a��|\5u=1���y8-My�2| �ڥ��� ��+��{��9�]�G�R��y�(,n��jfI�TQ�lF@/W�S�r��:+�&�;��^�)��y3����<�	�Rqx��ʅ�Tƾ�Nb���j�����ǀ} a�Բ&]�,)h�T�/^��v/wB����p�Z�S�	a�ې��]�$SY��k̀�t�a��}g��.�����J����%.p�-�E��Z�)��s��N߇P%��n���1<B�qO(�~�/_�%7����#�,��A�,t �����d�%%�v��-,+[�b�`!rx��F�`�K���9�q�G�\y	�ݍS )Ԋ}�c�B���o*�GsS��I�z�ȳ���&߫����"ܸ!g������?���e6C��8v�����LSd3��ΐS]6����}�M6\	�͛og�X�g���fS0���[9��]�f��hZ�.�w�a�+�@-y�b��eXl��ƥ�t[�`��1�wĤ%>�OZ�>��]�Smѓ���d�g�؆��fݳ�ik��ͼx�L���t�`j��� iY�����R�Ϻ1'�j����n�������K�J�D�vL�O���ɵ$U��g�`%E�+g���6�"i���iD_|WW�UC�mY�/߁���$��ܓ��7�"�S͹F�O��џ���I��E��u���G�oOC�r�醡I�/ >?��$�B���Аz|�ݤ�X�c�&D"^
�WW/�:����O�+��gl~[uB�c���C�\������q���o��bZW/��p��(�Q�ꋾ�)i�y�=sdeg�� (P��ć�&�:#��i#���pTs���P�=���8�+&�(�۰��������-�*~��C��Wv����	����K�����[�y�㾊�ba����E���j��Fǝ���cg��y�*3!�;�k\5���j]?䤞�P&���ݹo�d�!�|�������WW[�(��1�a2'��H�F8f�/���gC�{������Dn��Z)�J���*47��l�����Zt�XY�0����i�B���O\\�H�j3 ���e��]�ԮKۜ��F�"K�o�_N�CiXf�Z;߃|A��˯k���lQ�f~�,�G"A��-����w?z0�Po�����N����c�}W��j �P�׿A���?���+J�@B� �6��>��<�d��lR��?�ِ̙����@w4�E��Vsݚ�Vʥ�::'�)2��#OMT�M�{�Q��'��^�v)���3H�$�{�Luv���F��ʹ�5GjM�z��#o&;�$C�ם���x�7)&�d��e����Vs9�������Y
T?O���k������+�k;����0��Z����|��hu'���kٜm�����ce��`���U����7���C�= 4���MKDS��N��c[	q��,M����TPU��+"4������@l���.���kM9C���l��
��MWB�	�f��)R��zdA ����H�1�����X}�7ы�de�*<i�-DB!=�p ��F91��O}f#�zz�?M���Q�~f���Z8�N|���a�9�K�U��J*J��]%�WH��۾[�<i;;���Ԥ�e�N��]R���N�]�)�um)׊][�.;~���"_�׶[���Z딙
�#2u�qS���X&��5��֘�tI0�.�^&����7� A���;k�Hgv7�q	�<{����4YAŢ%����q��r��y���F�[��|Q��깸�up����ㆫ���o;��4(X�j���B�`d��3�'ӥʥI��(�!��K�%�b�!3���
���ܸ|K���4,Ec���7�N�-�M�J�Mp�8��d����|�mn�'��ߜd�)�ů�l)9	/��Q�N=�f�n���}�:��9��Q�DD�o	�<Ky�c��UN}'?�*�y����W䢞S�yֵrn_6�7Ll�$a2�3�h��0�)�`��<$HeWK�1(�
>�4!&F_|T�Xh!BHzO	��zo_w�q#@X��g�V��x��9�ձH)�����>�)~����kVG� �)��D�-��9E:o5-�e?������z�,oeW�0���Y�;��A��\�S���@)3�-'h ?:�����p�P~�W�N��j6
i������z��HK#!ḮI��x�+O7��?�"����h&ϋm����簒�������ʨ���k��݃\�5@p���5���݃�����2��r�}�o�?XÜ�]{WuUC�d�%"hI�A���9��0л�^!��t��h�G���9�����H�C_|��"C�&�C7�١L�q�W�z�ԟ�ݥOS17����yFYLH	��U����HKg��,����r�~N`%l����13�V�n�h/�?��T��:+@M���Ј�~B�C\� s�d?�J�B�E'?99"}h�����
�KQ��t���R;�zp��z��zA2��s#��ӥo����1 �}����I���j2ռ���o�g"N$�����_��N��e��J�2N>aI��.��ŲA�G7$�e+�O�J�\�(@��˛P�[i�-%-�T�x����{h�������$�di���JMꈾ}��sf����:���V�}�D�.55�u�<1�U6�D)�2��?�W��S5���������nm��/d's�Hþ���*U(ΪEv9�������խ
�����|�Qb��u��P3��o ���4s�ƃ�����J���M��=8S�h�����X��}��alp.`ǳu����ؐ$6�M�J�::��铑u���+_���v�,�Y`��o�����ˠ��5uꝽâUÐ��(���������7��#
���\D>׷>�9fQ8���P�.8��畿������� s�.6�c�O��UrA��JAH�byn�������y��E�J f!9� ݌�w�&X�?]��X�T�;d"�L$��e�TI���
�9��O��++c�yHv�<�2m��5�(FڧQ�9�����"��w�1u1h��o�gU���k�В���]M����'G����JƊ��i@
�eBo&���Ȣ�=�۩J�]��k��g��^s��pͭw^�P��F'�+7d�ɭ�|3|��I^�Lgm�{���ͺ��*� Q&7��Q�p
���mBYj�<z��o���D��EQ��[�jH�쌙�B����T�%���蹴𵿡h�8�tOr�{onP�QBM8���z���-��x7!7p?�}Ib	$�<�ߣ𮃂�3&3w�S$�/�'�Υ��+���40�s�uh�hl����!~ޚ�M�3@F¼e)_��m'q�57/��t�W��N�2�I��r����e|-����NP��B���Z���o@<P�""N��F!f�<�M%��ј	4��kA��?R}}L!�9~��d��rkw��x<�,�N���ᦖ*M����b$�4&leN�ߒ�Da��a�C���P�;�h(턩(6��(%�s8eD\��v�b)���@���8rA74��EށH�V��dnل|˪����I�l�dt����`2�lq���>q�	�|Xe%	,R�EbV*j��6)��E�R6��3�*7D�v��o1� �-!#��2�Sp�5D���#��"�����w%S�8L9���Q;��s0 �\D�Ѵ��Ҁ��s3��N.y�l��V�8�hO멤���=z���[��N3(��g�ׂ9�5�:6�/�F2o�}~�r�.��K3�Y,�G�����6Ũ�<}����5�\U���	~�y�������:"�'g��}���x>��Ţ��)4�?۸_d���
����;��2Rx�ޟ����}�sJ�=�D{�o�&�����>��%"NQ�wܟ.�n���gӷ�o.	��Ix�<q�$X�񻿔|)�@��r�\y=\�e:�p�G0�=�ܯ�@�����{�y�C�$A��h������>v-�G6^�_2`Z�b���*g��\������)�+z5�/>韏ta]�ekK�)�M��Up����;��*��a���Rxx�-߳�.�ESXƊ�_��Z٬Ս���+߹Ҁ�K$��`2k�Or!��4쓗�l햿���Eei]���L�!����͋�H,P���mX۬���9.��cIp�|%k�&�8Z
m�Fj=Yj�<��ꗦ�+�k�%@ΝBi�MI��Ƀٔ����02���v{~�����U��i�YF�E>��G�6�6<�~gɸ6Ŋ"�l~*�_keNO�ӷ-':X_P ���Go6�s���ښ�|������c2kn\Qn���|Ɨ����)��A����On�!1	̜Bܙ�Q�y�m��Vec"�u�6<�Ot�D�WWT@����U��)�q�q��1%�K5X������D�bW*+�5�C�&z0�����O0�R�	tȁbF�N����90�f����y���6�O��_�"f�Ug�u!�>N�؟�ބf��l`@�b�Ԯ�6�փ�$�)���?��5�����������QZ��KM�j�N��4Q���	�1Pf/�8}��ٲ�el�@��=���qr!����܀���2Q?2��xO���o��߳�����^r��)1JU=]B�����	�'Z(��P�LF{�� @4gǎ2&��mV���V��!�|4mc��f(��Ad�|z�ׯ�3��C^���S�2�Ѐx����.�$�����Ѧ'��b��7�	����6$���ƭ�ĭ�b���5U�`
7��(�}���E[����r��k%��F����: ��>��N��O�Φ��)�uS�w^ju��˨b�B���D��\\�+)�C�G�a<s�l��L͎M�;4���OU�CyL�Oc��� �c�����I��WE �O��N(�-k��L4e����d��ř���tM�x������ԂR߫�`ak��(D��=��q7��i󥟨mFA?��7��V��V����#HP�֞մ��X�=��*��$\��U���&��ˣV�n�]͛ނF�6��__L���cS�ݴ���-��>������!�Qrl6QY>��I.��!�$�Ĝ������YL�uU��36z�e�6��,+RP@W��˷ �MHz24���x��I`� m]�0qa�s�dzd���s�����)���*)n���������\��]M8�B~U� �D�o��u�����k�1�5�4�bL_.�|���w���[�W�N6h�`��Xֹ0�D�h���?j���l�.�ꚇ9kSQg�n�y
��D��ײ��p��&��k��܍�ޜ�h���Wf����S�)'��_��@�|S*��;mcyg<^����
v|<��=zW�۝�h�Z�j�b:c ��O��D݃$@�R�~$�y�"�j�~�+�������7mj$��q�d�V2l�ZHsrr���d�|�5�dp���܍�ZV��]mx��pP��G�ѧ�-�ׅ��q�W\U�]��f��}���2��e;��H�b�����O����.uȹr�=�j�C�? -�X��E�)s�!+�ގ�0� ~����a��%	�&��I_OA�?}�a�GKk�pw��4x͡�������s[S�Ղ��\�8q>�X"�D�5Ɍ[ke�C���s!�47m6T���d���Aސ�[PYv�x�R��L���v8�x���-���� �%�^�+�c�-*Q��(~����nI%����ͅ.<���:����w'�� q�$���!������������כI�����G�C>�/���6<��֛j~��c�<
�sR`��s>u��*%�'-;H��G����*[\'Z�	��aO������+�B�$~��]n\�J����4��9UT���L}�D�v��[��D�5���6adY�W��X)< FY+���ڭ�v�Ӌ���!:3٤���G�T��{+B[#JPuuwߺ�lit�'�z�wb����.�nAc�@7Ӛ��2�a�3�8��Ko�e'��V�_��t����2$��$��hgوLъ����VRjP�&���<�࣮�%��zl߾+�-���B���-@j��ᕫ�x�V��q�g���9/p��u��,	�P��p<X<'T���*�.�a��~llL�Ŏ���r�#�.��+AÄH֬�=��h{J���$�S��?�;TjѦG�uғ���K��ެ���Y�!L��QeA_�`,�v�\���f0�Շ�-4j�B�o��\�:x��x���qJHX*�2ˑ
|��֞X�*'·��ܿ�����	S��v��bW������=�[��#��n@�odz��8X����W���R2Y��vV�cn/_vO������?���_�Y}<���AT�^pwI�k�g<<�ƹ|�W����_.Ԁù���'��DaS>Z�g��K6Ӷ�цE�_��5�y� T���꿕r3�O
`Y[�FX��6>��K(:�.���M'��#s�A0v\�$�;��E6��龈����-����[�����_}�h[#��DoB�X���It���=r��v�݂��I��9����U�Z<w���Ӡ�*���V��dy��L��&��N �P��xQ�����FF�V��ib(�z�h҂X�򼙎��-�SER��mQ�(�#e��Ø���'Ə���^�D��jYnG��K��伫����u�ᾫtvv�`�>��B�'^xxXۿ�A�ـ�t���+�Q�Ј�2�W�eэX�S��6�Bw�DӋ3N`���2��ԑ�O�=9	�Z:
�po���mF�|3�J�����m"6�l6��4Y^��Q�.��KKѫ�Pb����;l�in6H�l����i<��5y�>��V[��0�+MI:^f/�
����`qn��!����6��I;�^-b(�N�|:�ȒY��}�U�SJ��n#��s���e�Dˊ�ݷ=��C�2��O.�(p0�i�?�f+Y��"�Ç"�-<��,������=�<��Փb��'*}�ɨ%���\�Ʃѕ7=����f�7Kma���`P1�����-וҟ��l�����iu��-M�x\����ސ.��;q����,&]�N�����������=H�-!s��a!��q�Lv	u�����ѱ�~י |���
Ӎ�q� �5ZAk�ªd\+mJ�\�:7� ���M6s����Yj:$5́����
��o$����P	��݀ƳU��8���_���,L0���:a������h/m��eg��dn{�� �֛a�(��(������tM��ɑ�W9Csg�_�W����8�L��1��*��q�i�]�1ﹾGU�@UV�H!��Ǟ�f17l5�\���rf=�II�P	���s���X����8+�(Ŭ��>+m�W_��0,ed��Xtv��:VD�d���{�7������h�S6PQ�[��0G�K�W(U�!��V��&��r�gO[-�D+L��*����~kD���"�j�2�]W�wd鿻�v�sZ!C�u~�^�U��h�ԙQ��� �:��x�k����(ޚ��dw�ѥG��{�����&��t�Bn	��z�K��pyZf�> ��ђ�)�u8G��i�׼ #��A6Q>
~�k�V�i�'�Ȏ�3��!P��'D1'#�}��[/~ɟ�ƃ�	+l�t����t��ʔ٨�hz�MLD>�˦O�T���[opi�W��|,���]I ��H�u�\v>�J\b�	��n�Ã���P'�Z�wk�Zck����|�%�����ߕ% /�ۑ��q�_���$3i�W��+���O��2ڡV�����/�~*�&����[�#�0�WD��-�L���4�?�����.�xKi�l<Bx� �,en6�չj�px�>_���G�0J�0\�ֺ�Q�BO��a��~i���^����[x�����s�՝�l��6 `J0o�Ұ�B����I iج�D�C"kqiɘ��t=#-EvO �W�����̟��*|��͍����y����@0E�E�Q{���F�������V�w�A������A}������������߀;rd(��' <�=�3��Q)E,Mp�#�U��p��O���F�#�$�/]��уg�M������$?lK� u�R3.��h���-N^�%����$a�h2O�k0l�/`�A�I�^�F�3#d�-ۦIׁ��t�L�<�$����	i%�g}��p\�T�Xq������y̛	�z���K3��-ō�j���~\p<(�Y���"�ň����
�~�-���J.���Qa:�$�}�U/@?B�%"Pt[{}g�{qvW'+#Y!M�	ײ��B�n�H��m�[�֪LRD�dF<�e��݃��ņ�+Ju���/�&�QL3m�C��ƴE�b�̡W�w��)]6�۽7vB��-9��4k���}���/G����|\�] �F/"ȋ�*�����F����D�а<达�,�l�7�Ѯ�m��_�ץ(��)h�y�j�|��'��&nO1j-����/���n>m�F6�����?w��}��q�Ym(����!8`�w�-J�6}�-f�Ҝ�.����v���a�qzB���9^����ٟT�N����$'H�����}���N�"�/�u7SS��O�6�� � ����@�D��͹eߘ�y򃘨���~����_Lz�N�ћJ�A��j�hպz4G�n:�6���:j;Iُ�3W�B~��",�<�TL^��s�!$�!��d��@�e�w�~������	�|��lX�Ӱ�*�e|_Y��ѩe*���#��]�$r���+���kr�/Lg����v����Ikc�ՎhÈX*6_�B6�[��Ƿ/��&|�p�T� �LRQq,��Vm������H���f�%H�&Q7/@ߢ?��X�w���j-@�UCc�*�"K�*�&�+#(z-�0�Ϣѐ�|�GD�ՕhA�7��91a��3_��O���[	����>6p�1F�z��R���5��Я�I��Q0$�d���}�x(>�}��
�:�3���A���c):��ۡ�x��N��>��KȲ����~�K��[����m����z���� �*"�.�w0K�K�u����t�ZI��R�������F�|B	V��'�������x��NV�
�g����o�������l<8����œ�bx��{������������O6V�����MA��ϡ������H�ez�~Wc���a�����d,a��)8򩱂�Cc �7��Ǫ�B�?6ː+Z����� ^��� ���+Q���g�p���$w�u�M{�"�eӚːP/�^�A��^u���3X��q���^#1yyTz�����1t��^����#�������'�d��q^I�j��xo� �	����G�S���=/���9ຼ��ܟ<�[/^��_�8��*q��jI������v�5Sk`��Yzj���&Fk�	��������.����F	=�_��g./������g� ����B:ҡ5Y��0n����F�a8f��ht�'��)�Or2K�ۧl�`�d*���3]�	ٮ�ւ��� ��[|VM�D&�Ƃ�nJ���>����@X��au�/@EHHK3�����`��7s�H��Beq�_�15�\������i��he���};��=J�N�Z�ʪ��ɛ�%T�3��*���##r)������q��{��g����� Z{%�п���$�%����F��إ�ր�`O[�r��GFmsS`��K�!0�0i=x��o��"R�c�il6��^c��Ul��"a��;n�q�`2sc�I4)}�����B�Z|Bu��It�K͟�ۜ^��Mu����t�:/kl9��pJ4�����.���%�������"R������8Q�n;c� ��1
I8���V�,Y=��reay���ehxﷷ�~9�׫��//�`��]'�Х��]���7�aMȧ��ScN��ܑ��qh_�����K�/��A�J+^0LRБ��*�$��(,T7Y'VRK\���>*�@޼�����p�u��]�!�w�����2��3HKg�蜁z��})�r��رRB�zXp�5���;C���Z�F����w�J5��Y	 ����"G��|� ʨR�Q�t�2��� _��!7G��+ L�H���kn���a����bG���]������8���mKˆ��Q��Y��:�h
[T޶��w:o��S!L����"
T�Gh��#�����/���x5\�#e��G�~D�r|�8����0�]�TL?=��+��*
;�	���U���c]',�����&[FLU��A����p��~�5�
e�mԿ�tū�w��z�_�?w�q~��Ԗ7c0=#�����3nIF<�L�)Z �wR]��2p�臭!�t ݹ���b��	��'�(Џ�`i�3��\{z��÷7�Qx�❥!�K���x�b4)[�������f�"�z-wy��c)�0�KWU*���9ؖ�خ�.䪊t�������6�BuL�%���
����q`(j�M
��{���?�ǲA��.�J�|'�����z0/Iꉜ����x���������MЅ,^��?cY/��m�k�	}���JPa,!��3��+��>�3�W�i�`
&M��68<@�TH���<�,-/��������L�3\y�2qn|4� ���?�tv�f��'b%���<�ڌ(��i�MT��BD���B̂`���HU>���s!���ȣs���&I�n�E`�E J���L]���ٝL���f�>�>0��jʿhw�'3���"n��(�����?.;�����*������*Z�<�	^��m�֙㤤�Ӓa`"������7�?3����#pd:Y`��$�~DEE-���ӧ�jPC�\�2=r��b:W���[o�P|��_ʜ� �������r��b���9�#Q��k��ž2���f���V��!�g�';�B�6	�k�$V����gh�=�M}�M&��m2t8��-K��k�x�7��������)�Q�n��)�I���pe^���<��G���7�K�q�c���ŸN��"ziE�� *�������P/���w&�?2�ޘ�ihj�'�\�C(0>4�$�(����* [�Y�Q�|4���UZ )��4��Q:\i'��#wv>7������F���#<�a$�,��ܸ�p��d����J�G�Z��`�� �?��mj�y�����ԁ*����
�X�����[� )WW4$�__ K��0���W�OP;?�5LM�|�r�����lp���4u\�zCA�J@���h](0�[�i�Y��\�iō�pT=�B^^^?���k��ۏc��~t�ɹ�Y(K4ʘ��פ;�Q�kf�.}���2�-ދ�~���^w�����&�io$���*�S�g-vn�}mmm���Υ�v�p������GbC�U�M9�K��R���)ګQ#�`���FЏ�Uj&���c/�'���n�c��֝Wt^�!��	{�����p���,]���c�5�n+��P���G������U66�¹[�ڵmt�lF���fU ~�0�^�;�455�*yS�VQ���@������ )�ڹ��-kO7]Oz8^�6ݍp{Hb���k����D�����["����e���7z"��G��n�h�*[��� 㰙e�(@J]iw��;sG�ǚ1=u(F�%mU��М�F'L��=�c ��NR�a���l'�жl�ݿ��ME�#9m���B�����Sh�la�<���MﱪN�.���B�w�Zb%�3[��0���zg������QgK6)�D�����,�ʚmM�i�y�����pJ���.���3���:h�����#Zܦ���7	|���+M�g�\�	�?m��|���O�7cO��+�P�F\��p�6Gea�@S
-5f&�2&�j��u�e����=-N����Mi�D�MϬ������r� �@ (C���Q�]��\Բ�5�{;'#)���I��	x ��9 �_==�*��ʍ��lV�Q��A�H��>��@5,��+��	������Y���2#�U
���g��ߏ��U?���i��n�8��1�9�ZYBԲ�(����Un�c�$�;ra$f�^^\�"�X�M)Љ�֙dt��L��Cn=>'�����yjZIZuK���JH�U.A��	sW��+���5x�I��I�T2{8} Zk�6���6�Ȍ�U*N�v>_�UP��HKQ�`eQnm��/�Sv�JUl~��)������D�uryk�'�@d��~��ÁFiN��������;���D[1L��<�?e�ލY�V��ȉ��\e*<���r�UC僟,�(��{3��4�E#��������JNI�ź����<l��u8��3��y�{�)1��E3�iF�Q����YI�y�~Oo$4�1�5&����շ��5I�K��/T��m���d��� +D1a��;�>�����o��7��o�%��!R襦JP88�~Ջ_%S%o�@���v�M���2�v_��_��ӫFh"��mت�7��t�̓F
��8ӷN�Eb�����F(}����fw���xN�?�J�����ƌ�y�Do��a�׃3Ԟ�t���B����oXyU�	�a"�]������bw����yܥ��in( ����`�-u��]��|{~���5��fD�V�^�w����*gǉ�DQ�E����f�����5e}��ߜ��9�4$m`c�I)���蠃7P1�q��ɚ��a#�N�\�X�
�"y����G��B���7��<��:�$�!	�_	��\cuq/�xq8v�Ü��M�d��%�>Q!u�&_�/��h������P5�*-�V�f��y�_�$�'�`r�s?�V�Ô��N�Rp<��ԃ����hs��#�@prM�j/�2����0D	����+�'��a��m�g¯�o��ʤ
�ѭ�F�B$�[�aHBH}�����T^��"F�P���7���[�w�=�l4P�AV#;v�N0%;y�S9IO�K��+1m�C���;���ի�%j.�򮉣|�g'�u��<��j�}1��]�)v�UK���S�L���c��$~��pc�f��)�l���c}�@E&OS��s�������b���e�D��E¾~�^-�9C�cچ*��ET`�>��"�UÛ��J�'�k�*G>?-���a+&z|�k�N�Rh^�-[��y��ކ�:88���y�{6z	��j��e�O�S Կ�������á(��b����9tN��'�o�Ǖ�����,I��l'�#d8]_�ɀYK"V
�)}��jH��Xi��	^2�8fҰ���f?���j�T g��ı��a�p��8'�h->�ϵ)��gm�-[����ӊxf��Oǃ&�jOŽ��t�$��m3�8"��?�[�}/
�;V��<�'-��>y���w���:v�ѵV�����8У/?yu�Ō:~�d����,��?����r7��,Nff������g�e�Z���#S'Gk��"�z��R�By�&�ed�Bd�d�$�dǵe}�]1	��HK#hli	����N	��ޣ�~0��s�c�����϶G8��I7�``=��탑�αS�:�����\�r�Ƭ<���-�p�����z�y��9����ak�}���S��@��hTy�ε�:��b����ϖ�+����Q!����Bޏ� ����M��$D��$�}M�6乆���g���(�#��T�z!s��d b��A�Oq�H6���S���$�E�������Yo�H��irA
G<�٢�&��L<Y����c?���P�k��s�0'Ǟbd��;����~ck�*�u>�:m�:��n�L��
���Y/k�z�*D4����ޝ��y'�nsd�?���_>��?�"���2��m�$ikz�ъ���T4ge,�W��/�G�O��V������o�G�#'^�./�g5Ho��}�^�s��>i��
�9��r�(�
ߘ�{Cp$�g�cP�iⅿ�F�b����$p��н�?��#:=��a��-�D],	�hu5Ɔ�MyRm��+�l>ǂ�+���-����~�+A��y�d���F���Y;�B�

�b5���Bذk�J-۷����ת`Z��F�_^hq��Ic��v|�h ��g���M3}v�i ڑ�u�p]��ӎ�O�Kϰ�'k�D���X�+`�:���d4�9�q.*d��`���f?�>X����+CB6)
W|*>ij���~��U�pޛC�ؼ�F�y89���t��gM��� �l�$�8��S4�~C<B��XpO���ZlJ���_,y�J�+)��A)���T7�9���U�A��a(�@5�j��ȫ/P%n&"�O�8=���ɬO��5`,&���e=��T��T���r�λ̱�=-��\�L��F2���0��/��F�+�L�^��9"���T�o���ra��hG�~��l ��/M\�o�2�z��PVE�w��)���*�}c.#n��mPe��ؠN�JL�kkdi:x�F0�'`I�Qc}��c�AB��ǉ-A�������Q��I����XN�Z�b�� 	�_�2Ǭ�n`��S��L��#t�/�mē�{y��s���+^�G��oB��m�}H��ף91�6�ʲ�-Y����ְ�J�[l�q�⫹���̔!_O�a`X�;w��;cZsx^{ބ��7��:�~�9�"Œ��w��:�������g�l��"t���+�w?��>_[�����<��z�=��|4l&F��gL���y�[��ȴ���[���*��f\.��gs֙*�t,[|j���"�e�[%i�D}O6q�z.]���_;��˰���?_�R�#���yr��g�&rЋGW��K|�S�~���d�a�.?�@G�׌�Y�����w�(����q�����̝���q��+��F�e-�$ B?p�vZ�,��Cz��l��t�q��缧�^��qN0��Q��B;��#�X��:�F���m5oW���C���X��W h僨ۑ�FY�V�iUyo���8;\��7�Garܫd,�*�wX�?���@<��iظ��9���lSM��vw���Mz��:����,��;�.�Ci�c��	��'��M)�v�zr^���6���S�1���0]��OW��(]��^%�i>�ʑ���������>Z^m�x�֕�����������K��J猊��P\���O#�uQ�oO�t�n�zu(��\�E����k���.ϥm\����3B�7�9YSLXN�{~Z�� I�������>�f���ȵ�gU�i�
)c�$v�fet!���3Y�rў\�ZU�.���b���/CUF<�x�\[�v�W�:/327-�P`R�^��e 6���Ν��_���=jC��S��K�o~�>�]������J�lf��w��֐�,�A������q淵�i����;��@{z��!�0�}n�P�2¤`-�o}�I;���(�ʍ�m����@9����XG�����ǘ:{�hU@�u�����=��ݐDP7!��d��������vuA̆��>:Cތ5u���ՄN\m��{<��Oع��U��������f�����b�]�&�$������g�̩r&��Q��'��ld˲�V�v�А�7�*�Y*�,qWK��nȑ�%�R���j�g�;w�d&
̇Q莶g�V6K��Ks��>��������Ǚ\K�E���P9j��|���-ڟ�V�����[�oٹ�ξ���.��	����������텘SQ0�a��J����k3��jiGy�&��'N>�Wm��/ჾ~���?ΜL�x&�4��1\
Dn���{/��r��R�<�P�Bl	��`�l�6���)��/N���EA�d.���b4i��Md�S�v�ׅ�ݔPyZ�M������7�
bE��)�xթ5�¿�vɐ 6�Ɂ�����!KwYt-Zp��L�<ۘ�/#]#���WH��n����k'�=pMu��H�����k�-��£��G�/�\j��+���B�'BNm��+��x~z�<Q����"�j���fn@�ŏ��XICxO�c�ƅ��e���а��G�'S䁆N��h����%���c=�Cb	�㽼#�X�䗶N�BE�ΏtYG-x��e��y��"��m����~����_����=Z���&uD�J���2%S�/f�R��*�x�Z�BUU5��SiN����y�R-��a�=��$����n̅�
�x��~}�]YPo*BǼq ���������j��w�����7�-����ٞ�͟��6k����4�K���:٘�?L���xB#�����Zn�G����rw^TXPaĳ��Zh�ĎW�5��Oί������l)s����^���"Q�D��. �	%m�	0PO)&�B>|����iK����C�����&;޲W�G��I.F�}��Xu5�w���ɓ�Y���|M�[,q'+��v����Ul�����*�~BrJ�����}Z
��Ѩm�Z���j\:�<�F5Y�^���9+�>���(٣a|�˾���BY�^7S�r������Ta��*��}�Zy��������b�L��u4�Z}��-���?u~CCJ!���a@0�\U3iF�w����3���F����Y͢�	�ʬs���T��뤅���Ikj�$M�i�?7ք��@J1[�+��� �S�!�Y���-�5Z[$z�Ěy!-�
�Wc�4 �Ε���=e���Ռ��C:��zm
��)MJ�юW���̻%��艇%j���BwQ/_���|ɛ>2�5���SH�(7W`K/�χ����8B�P�>�H����D�PUcl�E���_Ьt"����>�U)��������p�%��;��Qei��0��C�=���@q�qm���q5WI�;�}4�/�L�xB�(L�fH��[�� �肨�4P��M��xp�G����_�38��׎�u��3�,My��[���f�]6�\�-y17'��+��+�+�D3K�����{3I:x��+�$;q���wu,�c�k�}��$�
�R~���q�/"�/���Ԫ�E-�<=�z�v��@��P�Q^���^H�����:Fm-�;5,5<�
���7��J��fLD�_~�?�j��R
���8�����x������9w���w��H�_�����U����_�����S�L�Jng�ntY?sBC�}:��Cg����BD]��Bn�YT �����>�X�q����ո8����k$I~��˦�+f9�j�*�0.��ū�+����f����E�#��<]R�x�+|K�V����vz�t
����ϟ�����uw�0���)E���2���3����)(���"e��e��r<�4��Ȭ�~��S��!�������{�A�@z�@]�6L����c�̍T��weu���,dwE6�5_'P��zd����u/e�O���π5�M�K��`�M��Иw�zB����{ے{_>�Tf+����(�,L; �c/�\�CfMYT�I��b#��>���х���3ݑ�a~*�<�x~��sX��3������C���5��p�E��;����!DR=4Y�#G
�h����ߙ M�7n�������|����hr2�ܚ�Q��k��y�o��|@҂8͏���Б�>�ф�N��v��?ߔ(���W"��g'\��S���;��;;!=�o���4<g64A����'P;�Q�ᬌ�:U��"�6CAiau��P�ܫj\P�y����V��z��4+��5'P���������'�B�,�W��g��,�D�Æ��m��|׻����'"1� ��U?� �:>,tS��#�?�]�Zh��24��/k���l���l�Z���U}�\��yz#e{�n8 ��Mt�h��J�(Г>*c�9�������������)��_�x�5�1�WU��r >Dû��k*U��W/�U#��2��<��[M��Q�V��S�b	�@��	7`G/�}0vL�F��uv{�p܄�a��Va���^�Ɓ[���i����p��3N���� ) �:l��0@� uvvQPHq�HF�#N�����r���u�ƫ�.uUƙZmV��"Q`���Gn�G:�*UZ�a@�C�n�+?�AAYFfB��zF��1��Y=t>����bR:���%>>>G�XiY��$�>��Q�W0
'��̥��.6\�W�^��hA�Taaa��p-K�\������ۙ�-�����N�(�J�M�ې�������iu���C�6�b�y+�A��������Q�ZHE!�Eڬa��v.��P.+V7v-K�d��=j⁂��S�H�9?�wpϡ�������Y-n��((%��'�pŽI7vqQ���-x,��'2����M�'���	|p+���s��HIJQNQPߵ�guS��#ײ
�h����������D���&à%�(��@��@s�s�o�#�?6�e
$~�jk�2wlO��`���/�F���/7����!)/Q��i�95(�0�:\x�>�[�aJ�"M�q�'����e;w�G"��OԚ�8j�.#G�3CsĪ(��v-o�Fhpu�8-��@�>:�T��ͶV��kR���y$#3�)`�Z����������0�9�J�B�ì$I[8��*�,"�3���$�68��wHiKJ��8L)�'���艾��le����Ib��A�3���Xk3�vqu�ծ���W&2� ���~ƀ��]7��_D�rg,x�붹7�V!�����+�m]Ro��oL�f�&.\�0q~��)i�'��A�ϴ��
�:��0?ƹ�ԵbHV&�+J�E˨�R��&���L�f���5����ޗ�˙�9Ca@h�Ž��`��r.3STW���ʪ�<�h�d�P�M���www��.��	���@p��$8� ����}��{��ڭ�
����r��+--۫���ʨ[�^C�ŉ�3a�R_�7I<jG|\)����� -�IW�)�k�(z,ؗ4v-�.�3@���OR�'�5�h
:S�$TS�M�]$]�1k#���~��f���S�y/>mY�Ke�cN�(�C�����]�"�kTi�,��g�O�ͥ:3y���S"̼�m��*�o�ˇ�1">�w\���٭lQ���y�1`�b�}�U�~O(�m���&��JR1j�����u��h*���q����:`!kIKW&�F�C<��Zз~��K�|�i`��ɡ���u�n8�b��Vӿg�Xq���]'��kj�j��@ۙ��y�a�kF���H��j����e���x�;&�1����p�u�{�T'�ux|;� �Pt����^�,q�p;M9qѳ����>~[y=�\��_��bp'ͦ%߃��_�������g��x �
:7���!�U����hў^�R��Z]n<���u���ܱ�"�D0b�4blW�1-��&��9.��J勰�c��֞d{̭�K(ZK��t#�GXi̳�]�Μ��v��;�b���
?U�>D�\���3�U���"phw?5�x2��+����|���a���>�k�|n��o���X7�E7��_�:D��ҤL����}*֎j�R!�E:�kM�OO��x�RϷ�^�f<y��f���?}`ɶ�$R�-�A��*�����������榼�/� �c�ަ/C=xCW���Kc�����(2�P��=ÄT&��{:�1�]�7u�ڭ��w�"��/�z����xY[��5���6��s��3�\G��k Dp#�J����{b;�?�2�[��L�c����S{|���dx�0o��7T����*�RB�kGM��ާ��~٭��*���]�j��8_�p��m�u«VR88h�H�?��e�vH �#�����אbu��,$��Ga̾�ǃ��D��*LD�Ijڧ4���r��5�ގ�/Q{��>�;���T�آT�T&nfF�;|qqau/,(�D���?_h1���K0#V�%�7�G�'��F�͵㨭���m��,� �Cs~C�{��zv�w��G��;z�3�6hL��σ��pa/�V���g��āH*�}� �,i�ow*b�����[�Z� ��u��.��F���u�i��$�5=������-���ݯ�U�G�#�	i&��,)oS��{�/������PmvG���7>�'?�5��D�G��uk@�F��o�q�<�o������/Mx" S�`ߨY:^'�Pm�#����.��ݢ� 	�
& ���J81�c��[��Z����'�v�����!��}��A&�yyee�FՉ.}����ߊ�oV;i�ܡ*ʪ7X��=��/����4�����$���G��bw�m�VԚ1��"��_��`�x�M�M%k���^;��������������'�!:)��t��$�,���Q\u�}�Qo�[����@m�$���zpK��-ӊ�4R8'}�I�	8T0Q��D#�t�j���YҎי[���^ڽxY�o&t�������$�c�u����`�&�\Owؾ7��F�j���l�P�I]�n����z7��Gρލ�?˟P��6r�^O>���b=��/C�b��_+;�����A��&���tU�؈���Aq4�P�����ǩ�ף��3�z~�@G���Omt1C��"����,�&^mGd� ��J�!�w�<[W��u��^J��sWI�|b�h5��:�����L���\?�5�)-U��##Er�����7�e����R7>��"!�۲�ݪ�����0g/~���`zmW�y��Tc�
K��>��o7���s|�01fŽ<~�z�}&Y�����
p��vZ�P�M�@dR��A��k�;�c6Y
m\�����Ꟑ��������T�pj{��p��	�|���u^_�E���
Bd9?�׃�齴����eo���{G�(��. ���h����b CY!��J'��:̨�E���g�>���W�
_���З����M����ʆ!%c&�["�e��8s���f/7˙�P�������)4q݄?_�i.�<��؞5����S�Z[���O�a�f꪿��%�G!}���֌M���5My��ԥ`<b��l���X/�xҺ��%�[�C�D�+P�?r+䥠�x~X�o�j��8rQw:w?�����uH�XJr�f�Lp����p�`�`6$'�o�y��R̊|jB�ip�؂���>i= E3�
B����	�`.�~�[i0�u�����ڏ�N�.M�jr�M��W	Xn~��~Ձ]�W�1�+A����z!H�;�-U|��˰����@��b��+n�M�,P�����1���\��R C_d{�X2�>��}llX�ӫ/v��F��¶.e̅]6����V���3�|����D�rm�D	��*$#��T$d�xހ��� ����c$2��^��m#�D&�?Z ����O����t�����E�;��s���ޮ���3����C��d�µ^Ml^=\�c	ݟ}�'B^��׺L0-�qA�ow�i�~�o:[8x�°�:[Ŀ��|��'��$i�����T�
4��7��U}8{�@�*]k �4��Xg_����]n�ˠ)��	.�(��R�����z �X㙯��=���*�2y��I�ur%��O;h��r�u�[��FAz�m���|�|a�%8��z�
�o�~�k�l���ߘf�0ڇ#�f�ڮ/G�ܞ&���HuHӫa��I��Ek������(��.�}U����{nu��A2�,-��p�����q�-������Q�2M����r�՘���":E��Pl�un��+�D�v6��@�u������zS�`,!���}�!�)8�������l��L�f��Ď�T���TЁ�'sKq<�Q�}�sTC%^:�Q��M���2~�\����v�*�|z����v�nnn������U���Ĩ"Ϭ0003k,�2�:==�h.KG�4��n�Ƨ��j��JMr�k/5eS�xi�#yY��7���60��#i�}p�mr��W&�K���Oq~���'�Оԉ���9�I�4kO3���Aa��k2>}��,~.�Y_�	��;�����u����Q�;\��|úD��g@�)̎!��ՍZP*�+��Nql�-��z��._<��S���v��Q-� �:�*�}p�� ����a�<����>4��D!�@{��Jz`W;�]M�`��f}c��6jy�mέ��߲���>3N{{;�jj��\��Y�A������+`�W.�>��E�0�3P�H�����rP���!y)x�A4��M��ޢ�����WL%�|"���������fW���0|$g?W�>�����H0�eK�����St�t{GY2ZשP`Ӫw#�Q��n���O�������Iז �(�	
���
05�� ���`!�����L9o���3�6ஶ�7"{�UD8{x��d�8AU��˗�n�����f����'7w�6/����z5����kiǝ�,l�H3=▄@xF��z���\������" i��6l$�����	/{Tܴ;�=�|vBG�,-�<��2)�?J*+�O������t�N��< �%m��x{���c:C�����ԿރJ=�.����%;�_Y-�n��E}f��4�fU��/�)�z����{~ ���es�2���p��^R�֖<���0�r��HS��V��g,z� �p4��N�^�N�`�`F�l��9�ЪuT�0Ԉ�y�[`γ�&M5�?�e��LCD/7��S��j4��WW���jS�@����}�2/���A��;��a(�s�K�FD���82��13�6���r%�ŀ��Ԩ�eҒm`=~�˓Px�����F���U��5k�f��F���BI˲c�>��Гy{}o����|�2�!{E��6@�3I�����H�4p5�N
��ǘU��ڠ���
�ά�#2�'%�jmN$�,�^�1�z̸N��HH�8���� ?*�V\c`��bUw��}�ȵ���Wf��|�I4.]��
��a#F���;"��j���:�䄜m�N�ߡ�P���NbT��;i�j�r{Xg��"y但�b��:=��dµ�?-DS�+��3��͡f����e�A�29Q��q}pi�N�Q�yk��P��(ԹP��D�^^�ۺ�H�������Psu��?v�g��\q�a���]�i^ E^�����)��Vi,������8Ͽ�jT=p�0�]cl��ө �x���ͽ���c�*��G@U����J��_ücx^��DQ�v�Qk�LA���D"��,=��
�����Xq�Oc�)�q��i���6�����ӑ��J���8Fd�x��0����+���id�.`ʌ~P%���P�ie H�C��h��u�[���ͥ�"��Ks�Y<��"(B�	�:�����.�!F���H%N9B�;���\�#V�-�5��$���B���Oc�z�J��~�18���2�3�Հ����sj�5��7���-ړ�FA����E���W[=*�|�_�#33��a��n��d����>�N����9\(ĭ��F.�7t�5�6!
�
`znd���{��?�bT�������K?ီt�;��J�H��7^;�i�M7 @����8<�:�"�x�v��$2�Mӫ��D��M���4�hP7~'�Y9 �i�(S��ٛ�����'G8���!enme�M�b�ɫ�U&{���q�Q�;n�كf�x�mt"�6B�h�"�ڦNj��/⤆�˪K���b+Z���>E��]�p�?ʶ��`;��'�6}�n|8Sb���&���/#��eZ�{A�l!W����w�j�3�Z�����'�63�H�H��ys'ƧħRU��ճ�բ���~�3'֫�9�&1�1�#�>Lu�֩ki��)����CS��>�)�$�K���dq:�8�:� pdj���Ƭ��Ԩ�\�����F1_͌+����Ʀ�sC�q�eHY��b�� ��`����`�.P��7��h���'�&�Og����F�.i�X�S9�gvh�6�0#��"�ż��A�.�W9���{��X���<�u�1eǏ",+��ɉ��_�wl��j�ٛ	�w;'^�V�8,���8���-+�3��I�@뗉���`D��G"|��r��}&[lq��y!��kw�����5��?߶[�I#��5���\qVMd���\����yS�g��7�~s�mB���TyKZ3/���;��t��&���ᇭ�L����r��R1��3��Fr��<i+��ٽ��h��ӄ̜:��BJx��D��z����&��wY�����`�?%|��doC �hJ�|
:��b�U�dyݖ�]�*���a�'�!�ǧ�^���r����L.ۋy=�؇%Vx\�):��a6�;B��`�1�Ш@v>����.��ԢҀ�����Y�uE)��s՝�S0cV�~��$;�n���E�j�`�a�l�&�s�� $��a��%�����^X�XH���T��4e���6\��.Wвu;���{��wv��Ios-{���>���O�4к��h�膷�l���܀�/܁�e��݄U��w�P��L�%�v��^U�e�A*#�Z��*JkKvF�I��Ԇ�C�5���T� C�\�f��u"җ���:	�
�d%��u�"�g�N^`%حY!n&4�΄q�|�q��r��K'חI(���q�X��{qX��uK���&VV�c���ֶ��Kv�W�v�ӡ�x[�w��N�9Y؊�����4��S�b�2L��u	F���J�X���$��ڻ_�1���Lzg*�'K�j4r����c>Y�!�[Aީ�b�%Pgf�gHhi�c]��B�,d�"�hh�,�V5KS##b~�DS�C�&�1���-��9IeN��N�c�e2J#�.���h+��G�x�`{Kݚ���=9�.A��fC? TɄ�)\3t��Ӂ�r~��R�Y�a"�z���ΓOp���<�V�Mrl���J�<M��T���]�b��}?�onF�Չ��ځO��.hw�籗����Z��gC�>��x���UjQ����:�� ��qh�t����0	hMd�A��C�B�*J�8L���'d��q�!���;p1�P}��No3�;�2�z��a� �?]�����v�g|n`չ��/�_w�$�e��C�a'�]͈��0���QS��2f:H<��|��s��6�0�/ǥ�J��^��t�=B���{T�����M!��A?gu��m)�j�HS���٪���R	��VI����Zn�u�3�mHhp���~ ����`��������8$$��|jZ��I�f`��,Q�����`�����r�x���z�b"X��&?oQ�n�"X���9.!!����T�4N;�u�ȎJES�D��t<1,��[c5��3a<����LZv���@��>������)�P�D��)�w�L)� �N�5��5g$�S��:M�J���br�ɞ����#{���M@���=�o�� R48��ϙL�ϴF�yuS��	#�a���Ip�>z��fh����Q���h�>�	�	|6�]�m/Ff���L>�i	�簼"y�L����4kɲuꙗ\\#��WH�!cI@�3s�M�j����J{1i�������DJ�1�9mo��ǟ��3����=H�:���J�gj
����]p���@���Z��,��\4��q����]��X��!�"I}֖p����Sp�I� %J9�Wb��m���C)���K�f��1�$��R��9
^���t��eEM��?��N��+L4�~rշ�F������#�����Y}C��g�t��1�"�.[B0q�����{�'Ҳ�6��OT��;O��U��Ԛ���Tĝ .�0������S@`�9x�0~�S���㵸v��]�b
D�t�U���EEł���Z'}��D�ܰ�~���;A��5"Q"~�Y�Hޮ+��w���G 9���<�1�{_// �����pQ,EC`Z�/둌�d_��j���|�.���T9*[[i��G?a��f&i�1CG��sy�:�����aes36{Fu�����ĉ���jGD!3��{�+K�0uǏ ��jmH{�s�tX�`�����m�zh�Olux��O�Z����q�xϻ����W+��[��v����y����S�DYjhldT��3J�e�5��ϟՊ�~�	����q���J�Ǌ;u|s�$ͼ��}5���;f�LaX�6'����`�,/L-��V2��m���ki��w�8�>yk,N B�o�<��b�l܎N�s�<�_&�zb��q��4-$zQ�ݍ���c�lH�n��%�"_�iO��B�Ȭ�&�d7��1��gܳC��Tھ(W�5�}6�N�ӥ�ޚ3s�'g���H-���&L�����y���Zf���{%����j��"H�z��\[N��o��kI3�9��á���d7�p�sz���o�e���y�t���:3�(�W�-�l��^��aq%�{g���}�"�''�(��7� �)�Ca��ߵ���v�ew;��g�L��y�˩d�-�X��IYMHL��t��v�_��z
�D�H��(�S�r�zI,7��	TzJ�/t�	FB�C$ӕ�2J��]ڨ���ME9�ǽO�ˆ�*}��$��u�N��,~�ʕ����"�,Q��VT��u��Al��B����=�@�s<�=�����r���Y�1\0z��E�w�����n^W[E�����rDtV������^q����.;M��̿��8���w�J� ����։ߥ��r����=q��#exS�7�<"��O��C'�~D��]�<\!\����?��&�T���N[�>n�;��Jv�Pn�`a@#�@r3��x�E��Pl�״���!i䠡ϼ˴��7��$$�2��U���I	Q�O=�{2>��6Y4��)��1B����-6����=��π��.w�׮{�\���V��f[Q�μ�>�h��s���Bv�Ok��Q[�8��Ԫ1k�6#L�ω�Pu�b���yo[}K�c��W��u��J��A�2~U���qX��,//{x�/&�u��:}�z|�YFBϤ��`9�I���d�9?�}P�dtu��R*ha}���Ѥg��v�
S��p����K���C�ݕ�Ig�X�gZ�7j���5����氏�%ɏ�Kj��-j���'7Zsh��=��BX�[��	#Q��K/--�݆�9؆Z�Hb.Ó����k0�`��k �����g�yI����a�l�U�-N��q�]�����;e|)Ԋ�O|��d1��X�gbb_ ���%l~�T�-U�d�����4���Ӥ��6��']C���C�#�W�s�+F9��{z]�G��D�>�>#�c)I�uky.�����ڌ�9yO�r�O�t��xD���k*�v{�Q����5O#5	���/!��c�w~B�x�ŘL����vj�~�����+�U-ǩ��إ�	X�Y�1</�P�x��7�� �)	�/�������g����J�����V�������@BA1�x3�P�Ě��s�+P_�f�ˉ���dU
�Eغ�7�A׮?�?\/�7�i1�0��>VN�L�+T-^���	>��0깎A��ǝ��|�uv��p`30N�Znv���r^�z���:���i����N�Wx#��<����0��f�T,G��!�t�~6��fB[�/$�}B��!�a�YP��3�@�v�s�Ȟ�5z�����*���&l�>k�8�-��^ֿd�lA $ʘ��&�|�yg[�N�K��h؉˳���m���̭��Af�a����j*Vt}%�\���'J�=q�'ԙ!��H��<v��I���V~���'��T��⨍�%���1ڐ�J1Y�}Zƞ)A��݋��2X�7�jǪ�j!�{��1۾�<��eoU&
82
u�	��WWq~\"�3Մ��C�>��`��bKN;X����=Z�JT��a�1���TH��]��F���D9?_�=D��ՌxA\$��Y����T�BH��(h�)w��w��A��6�8@��J��3���S��g���&A�y̫5�o9l���ݎ�����Gh��6ټ�?�+^홝�i�(�c����y�~#S�No<��n1ꛥc�e0��2 ��r��ׅd�[�u��%����}��e���>���2�^*�D�X�	K���N8��6��D���������E���N������I:����0b��3b�cВ���ē�N��S�����7��	�D�U��9�Ԧ���0\N|Ba�@��@���F�3B
�)�{z�t(�P�K|�W�җ�����,D����S0)�C9��^�7E0��b�ȋ�q�^K�L�i��v�i��m,Ѷꀃ�:���P0�0p��u�wǍKU�󢢧��#j���5 ��g��Lq0Qؙ�G�cQ�_�37�<@3�������O�cI��Jj�9��\;RTk p�3#��#�/�RmF�

�{� ��]�[p�p^B1��ST�̢éÄJ�w~N�4:z�DhZ�1��2�̷�E��9;aR���v,�R��0�f4WD]�Y���n$q<�� .�����殷��w
�'���1��v8�O���j���N!�f1M����}��Us���f��.��]�'6��+W�}�Uf���ˋ�7�C`�e��X�����P�ۚ�������M���~�̔f�bu�b�DV�8�b��mJA�]o4�6b�6	�'���4u������t � =4����!��vtc�{�*��S����\��KL<!�d%�q>��x�1z�Zay'@���J�1��.�Ic+����?v߷����=�6>�C9���Q5�;�.l��N�O�/�w^���@ϗ(���*~|9	���.���s���u�v����T���1W��C����� u�2�z,hj�!n����s嗭���?�g0pB��c�W�LS|�%���@��R�]s(V��.����lºũ��g��U�u�/���e�C��]��d�;9�l�@���ZC�s�/@����Ⱥ�.-�hhu��]fn�<l��)���O������YS�WοJz7{�����<��}� �!���d���ۗ=�fNNN��mp@��^e�z3��������������zŏ������S��c0P<�\�����B�e�o�7Q�B��"�����Bv�*f�{�\?����ӔOz0��0����q;jo�O��J_�o{�T+�h(����w�Ȱj�*���RR:�C�7�gB]��в��\B����z�*P�0d���=5�Wk���R��ɇ>JЌ<H�w��:d�.��w��MLL����㿷�+�i�Ŋv1��,x=�D��������{�}��0S���7�[�*���.������س�*9O�T���{Տ�;x�N�\n鞋J����}��+w�3F7��\[�;�'(�I�!���(����W(�%��E�2�bC��!L.Wl�"^W��c	��z�s�ڤ����t�	uf�~|,�|@���|��a}ݯ�)�mv���R�/�%�%�mmC�A�*��v���8��:�|	�n��L���߭��q��V�z���*��X����ByfM�wE��ܑq���/M�G{�1�@k�82��ȕ�V��EB�5v �u��HE�PhY��8�����H����J�eʕ"�׷ح���#�oO�� ������pqڝ¥������e���+\��f&� k��=��|0ZQ�0��Ɗ<b.���1_�j1�u�oX��v�y3Km�S�k�;$��O�(�qm�7&o�ӿa�@F�vC�<�!���
3�q�Z}�v�%��Z,;��v��4�S�zz��~4�h4<��!�o�G�ݏy~ި�&!�z�4.��YG�e�2�(W��\ M�Sv�N��6�K�_�/Ow8�;��y8Mh�l�7y��-&M<b�Ol��K3��gr��,��V;�G���
.�W^��?���`�b��q�$�ψ���?NBW `�/g�5�̹��qj�R5��r-��[Q���W=�b+}G���'ֹ�~\ ��I\!L��yd~o������:#\�X�Tє��gm���O� >A����ʺ�
 ]IM>u�������[uPLAOm�K���'�YOdB٧�RHF1��9�;��Փh���|_�<=�6��1[q>�m;���`�y�g[�y�c�F����}=>�c�v6ɯ���Do�VeJk�u�3�祆��������N\vb�km�C���%���6�%=�˶���Y����:@�'�B�r��D�I�x(#��v��fʊ�q��}���)ֽˑ��N�����S�К~�,�?�5��B�l*��#<{u��lqs�/�����"7���3Cn�k(%��,��pl��g�19[;��'�@�E�j.rд�|D�׳�ҳ��C%�`�}Ԯ����$���N���7#��y�HSc�,�PE|�k��":GL�o�-�gg��������#��/���})�_��$�?��������prh'?��:���Ct�;�i���1uր��$�j���Oi�{6�q����䎷E�[ǐ`�u#���J�7	HK�&�s��2K��y�mN$�>��v�R"�u��G8�����Ƿ?�3]�[0���N�:�����h�
�;����]�#�������� K����E^�W����`-k>ܮ����b3]q��X]o�e�Mۄ)g��[a��D+@5l�s|��?o3�'W���t^ڡ����M���T�S,��0��DBH8�{��HJj3.�>�tq�~LH��Ҝ�tN,�!`n�\N�Uۚ?->61�C`#�ք 4{)!/S�
(�{'�!r�CF�bBh����_n@l�U$ON�c4�� ��	���3|]���lI"��
��EyA	�`r;Y����������Rl2(`K��l>`6w1�[��L	���.�7�syqd�3f���DMH�*w��C�R��^#�L��*tA��x��l�ȷ9��9�Lc\�����h��S���Z�L�/�9X
w�I[�k��]��_�9I��&��Whw���Jaܞ�޾y�o~J�&�9���0gQ�'KQ?M����7�q����񲦁���d��2����h"y�:��=�ȵ�_� �j�`��V��^��Ϟ_m�W�u�i��:��;{{�TT����x��S�+��k]��|:�e�c����KD����Y���~>h���VG�WD����sJ�^�*�!���21l����JX߆jp�]�VA�(C�>f�
5����C8�0n��)ֹ�VZ�0�N�����[�?N��_�څ����G�i���Q�6���4z���Py�N�p��K��.��$���^8zQ���<�i�7 ��₶E���)���xT����7?�ZB�U�+,��9�%��,�e�]|�&�҇<I)S�� 7^B8ۍ37���Ä����6`�b�T� � M�����C��io�b�3a��+*�&!���$I'R< \���� "u��Q�k�c�o�����g�GK�R�7k���|����Q��B�w��$�gɈ�͂�P�5|7Z��zU�o�~�CH�w�����jX�w�^5�8RY�U�3>ى�x����N-�������'L�4�e�.�Q����[�(d�~XiqD�-����"^i��j͑A�@��F�2��M'8z���	x��"#)�Mt=�+QW��ɕr��=��;X$��qx���f_��!u��]�4d�
��m�,p�u��y��|O���i2�[.k��'>h�^X��-�a	�8 ��O+/81��#���F@90B|��3=A��l����I�,ފ'�Yl��Gkk:9yy
!L�HT`��V�~���ҩG���WA��K��Mı��CK��+T�1�����G�"Ʀc���}������م�Om�zw���z�gB��
b�M,�RX7��O�ms�x@��O�w�k�q�� ]0m�������g����}^/T��0d��]�b'�HHz1�<�L��(TUUY�g(+]P9r� M�!	�jj�P#t:�̸�
s 1?��jĦ���T=����U�ߚD��|�jޘG�o|i����
�^��H�(2�xQ-�Pf?�?�Bn*˟ D�������.ܪ{��?7|2)��k�@Y�zB��<�~{��gF�ek�������� �OFjTkG���G⾻ �&O�1�3tѻ����]M��}x������&�s�����(B �>KHx׆wH
��g� ���bX'-)	G$�}X�&槮e �,M)ɏ�e�1.tz
������t�My|�¦���8ڇl�7�w�ߔ,v=pP��G��䅎䇋����d�0x8>�~�@l���2��heG9�µ� i��捄n�*w�!P`[�*%4��|�5t��t��)� Ȼ��(Gv�e��i�Y��E}����jٌ���K��nE�w�����Q>��ΨY������D��Z��qt������`Yw�iz��e�nc�~���ɣY���>	������O>�)�o�h(�b�yQ3�Ƞ��}�o�P��Y��#Q��XT��a�%1�h�f���~<H��~�í�"9n�rW�����y2�	�w���O9|g�l��a��]�c�/�*�1�N�0dXA����8�E���r�W!_nb����LT�Z.N��^c����>y�m��"�À��_���}̝{�~�R�{(K�Q�T~�?f��&~7�]S뎃~��]}�o��KFI)B�$D�F�Ɔw��n*�Ј1�煱���R �*�Ή���^���B����Re��T�}�y��T�<��I�'��Q�N,�6�G7�;p04��>�� Xj,qABnP�a�
���/��Z�wg�JH����a<b��񅰉3���q)�b�4|�jK�4�<�F����TU�)�e%pdSG�U*��%�חяN�Z�W�Y�A��A����e[o>���:�wڲN.����LhccSﺯ����ݕ7;�9yN����/�c7��6�?/�ˤ�W=�;Գ�^b�I:�K��������p�}�+�ѿ��y�E� �s��l5���q��+@��mFo�."�2鐳N��V�.�U�,�#R,�ZcSԺ2�-H�N�E�п�MH�HGG��w�v�=74UM��<�F�e����;��sUI���Ŷ��!
쏗[���i�l�67H������;k�r8ۉ�8�W�d���<�Nx.,���� �Ǯ��>���
T����^��]j�I�ֶ:�S���}{,ƃ��`�vZ��'G��S4ʙ�~_s�~�X֕������%����RmS�ȱ^�}V�\ q����v(� �P׉�>��ZӶ���⽟��zC��3B��'2B������yL��|>�������vr�Ծ�IJ��9~5k�_Ү�0�C��zq���~��M&�b�SZMU���+?E�ʹ0�g���1��N18�ˑ�m6���Y��Xn`)�'�ϫ��a��ֻ�"C{�1! x��PدZ�<��,N[%��㤘aY�8�a!2;� R���h|Q��D>��g���(�afz4����Fz�PR��4\y����lv�Y���%���y�YW(���	�K�*+/�8��-빐�ݴ^h��u���Ԧ�)�KQ
vYahTZ�����Vi�y���fB������*o1�hh�q��o�7������G�[p����<��e��7c�Il���;2��I_�����9<�l�Y����=u��EG�IZ�C�.�d��Z�;������VH+ڜ��Sq��w���K�R�~�0���-#?��r�#4ܱk.�qW�|�	�I��;���&����y���o����&L8�yx����	�4�F�������w��|�4����|Y�U!7]��ਜ਼Cp^q;# ��m��KUC@B�B=x�)�iYrs��kQ���iY6���m~ꇌ�^�z<oBd�����
��SMM��KF�AYCno�r%�p�e��CA�Ņ��niK���3H�,T���'��w�D9��m��o�3�/��	T�n�@^}F�c�cH��+�zk{+�i�D:��2��^�VM� �I:#�����B����#�����'߿c*��ik�{����k�s*�V����Ӹ~�5 6Ѓ� ����~x�i�:{��u�Ϋ��P3^��������e�� ��<��搋����y1`�*y��w)���~kL��S͛
5�-�p��LG}*� S�vw�y�������C(}�OLI��2<��	BO��P�Ol3Xq�a���� �n l{� 3�BPgw2z��n���)���b$B >��x�B(L�q���}ގ�Uz�MSay9-�x�4446.A8oV�`Φk���n��Oý^�����M�n�G]����r��Sw��РIq�oD��8��>���$3��YX� �7])��pę��J�eg���u�@��d��Y���~�n��g�o*��|g�.g���r_C�����#���F��5J�����W6'О�%��h>��pr������O4����P�;���m\�89Z(��!uS��F4T��/��}23ȝ'�W��Z��gw��n�s{��n ��o׶����|߮��\��{��������z!"��E���z����TwjX��
	v�d�]&9�yy,�<�*����w�Є���v`�0u�p��&�����-d�lfR
e�߸����-�o_;��۰�}��p�E�%����w-��DH��E)PY�n��\��+T�P�^���Z��@�5����7�p��-���{r��[L�G�!xvן�}
��O얗��n��}�y���l��J>�}T���lb�7h��!x~<�3<�e�[P[$�K{Q��wʈi𻉜����SXVzxBX�?U�L&6Y��w/E�ׯ�_y4�E&�������g.vi�k'
=�➜����aء�gA��{M�-�(�iwYӛmPQR�$�)ԛ3d�̓���ۥ��!�����®���_��8�f�gxYfY��P���9���7a�����c��8oDɠ29*+����|0���b�>-ܦ8��;C&7�V�~Bv}�&��r�Y�s��р��8>��ᵛ������X_CM0L@q>����{b#��cf4r�Wd���G;]'Q�@�.3�B�erW�@�B@�>�47,--6�ߠd�le0��I�px���`��6���е��B�S��y������\,��|��(��O�N�ϧ�N �
2�( /�y�U
�^������M��O���V�Љ���������@���B�l�(R/��~�)rT����O �z��JR.��l?)��-�a�� ����Xy��F�m�3_�G!T]���HOO��Ȩ��/�X�Bk����ZW�7Q�?o����m�FB!��R�]l��H;�	 �\�m�m3@h\�)-*�s�x�E�Z��-�!b��i}�I������J%�]o���E��ܧ���~$GG�[�q�/�o{��(��*o���h�bye��ȊQ1p���"ٳ��>�>Ze���"8WC��[GLJ~ߺ�S�ctc5��~!��m��jQ�O5
~����	�����-��!�-��`�5��.�5�ww(P�ݡ����
�J��`�R�����%���ͼ��@ �dw�������}>��Y��[�S�>k~H1X��v�3lo@�n�L���z��r������������0.t�>tu����	S���v�yH��m�L�?ߍ�� <�_\/WVB�� ��ܷ_3<��$r��Y�nPv�Ӓ��� ���^?��@��-�������w;Y=;����Mxv���]k�g�,�Ұe�@�H�b%��E����±w����*���Z����`θu�͒��ؘ��9�s׹��NP��O[���6"�8x�3���ź��zі���Z(�F�M��d�;J�;�*M��](k;�Q��k�i*�B�4N��O\����
AG�YP�J���7�I�{�_0-�#�{}��G*ԇV@��usG��mK�87F�YHm�q7�I?� s��4-ags(?ǵ-�𶢬L��By޾��;�3������յx��R%�Z?�.=qu�4r�2��a�x�(>����fj�2<,[VVf���a������y@�ލ"BVާ�(M�4\)������Ȭ/����\�f�ׅ"=�*�2Y�cB�c ,O����=�E���@�t�(�Ń��e�ɏv�!���TG��V��6���d���"t��!g{Yж�i-0�|��6�b�3i�l�Sp]S��,^�6�Z�:��A��v����o�'��c�+��'�������΂�##�
��CA�hg!���S������9*��Xe��q��
�R^^ͪ��<$V6>��¹�����Ȍ�:
x�*Ե����r�02��U*���񹸹A{�4�]����Г��ǈ��U�ϟI�n��E�EJ޽�F�����QL��欃)�(�ʷ=I,=��rJ�u�Q��>b��F��Y�W|�U���J
&*ss]_��*�|Ğ��R�ݤе1?|���t�r��7���h��z�I����#[�N�?Id׭�g�eZ������x���Ph�50�Fqٖ�$饚�_!��Z(*��$�ʂ�?���륶6�@#��TQFL}�{V���$�NGz��,�	�|H;�/�'p!�ch��j6NA�2���W�'�C����-ķ�P�M�X��O-����|��O��H�@�$��D���#��x󻐐�����,?���5�Ɩz���>�ўԇ�)���U��A_5��Shm,��7����gu|2��CW�������p_��^yѡqQ."����	]K�<��L.)y�΃�Կ�kbG�k�s6K��.y�A`?�����bG,���C�=���]`�� �d)-Ϋ�{���&$�*�����I�s��ӵ�9Z���
U�������y_C��Q̪�˔��(���/�7R�J8�uu����7yʘ�38�͸u{�V��L�������߬��8���@WR����.�k/��#��)��㫺����z^�4���<�Hx�9(aB�y�#�;O�s��䂣�<����I�� ����Ǡ/�-᤿3B����__���6��w���%ٓ�j0�O�	�Q���� �a^�21s@QW0��TT0\9_���Df���,Xu'?�Z��o[�k��J�d��@�v�5M��A��֖���6h?q�$�>���2f

����g�/��ް��i����3b [�縡�& �Ա:ztuT8���i ��!`$I��c��N#�:��=��Q��l-Y���y\4d}�:��O�+��9�<�G�=��fՠ�Ϯ��x�V��;����y�)!Sm�p959̓���$��� 
��i>Nv���;��u$��_�}���|Y�t`��<;�S��X�^O^��#[�r2�*謭�-G��m�kP[��f.�������,7/����p<$,h�T8qgӊ��UU#���-�N�sV����P7w���7����
42dif��ݾ��o+���A%�`��C��u6�|����B�����9o6��0{�F���ϴ;���V,y��5C���_�-��-鉾n>�BHCPS��P���e[7������4��G^����d���Y�o��XQ���le��Z=�����<�����5���;�,c�ρP�L.�:��kq"t������"-&�Oc�����v�˽����|�}{��ǭ��b��-�-XQ��I�e��:��Z-e�@�#�#q���+A����Kkk�L���<����
`����t}��(I�
i'�I���\ ��KX��	z|�lqz�K0-h��i!�������������ڲ����=�烽[)ƍk��UN��������(m.��+|&v��ui��bt��=�7k�y*�B�8��;�x��e��]��j�~�Vx�z�լ������D����\~,��_Qc;R~~��0x��V6=��4�F�(K���g3:th����w�n�]�Ǳ���F����z6�A�P��5��9�h�5mO���B(>cg]��B�S�!9�=#��5N�K����m?`��j"�
�"ϊ����e�jt�-x����u�vȾ��
����P����#^��{#*,���@_�>�鷘p��_cҥ�L�h��ޅ�8�*q;k��ҞV�F��4��;ќ����|=�����r�K����$tkI.��W��Atv=ojy}0�-�ö�+?��+~~��)	F<)�O4oߢp���G�wj� d]/+ʈMNG� Z�ޥ�1���|��UnV���~���w|��)��L��m6�(��'l�_�d8��Jg���"uy����3���GNw)d���n<L������)�3G�1�͓�z�J�Ů�uhBF���$����F�6+.5�g���F���a�/q��~��_L��y���&'	��u	{�<2��F�ڑL�R,D������+��H>_�m���o��8��C4�9�:�2v�7~q�GƋ8r&����� As���_�o��?�H�?Sav�&S�<���AD'
��5����ƹ/I�"u2

J�B9�a��`���ld9�&��$�42AL�.P̊�����h��l���l,�ur��{����$�p�A�h2'�g��6yq����� ���G���άfb~X!��	���DU7u�O��B����u/���8+~=�h��^�b���<�҉��i��-qPN��&�d�7�Z(�j�w����^c�P�2�I�OתD������$�][M^��_Ў���0��o�#���NP9��Ս�kN��ӛ�/8i��G0�Jc|T4{90L���*��~v$$w���~�$���Z��Mٻ��=ˇ���V
-&�8���.�����@�htP$
.���^Ye�uȾ�ߌ�{���/6jd�!bR�(F�>�aQ�wř߈�0��E�r�L��֙�H�X�a�����:?���0`��{C�#ӆ@[k�_���p�����h����L�M�,L�jupΡ�yi�H3�#gC�YqlZrsR��B���w�n"Z$;T�%���We���pJ��w�D��;1=�˨$��>a�s3�<}`#_�y<��E��5^p'��Ӗ�SAh�(əE�a��oی�q<�ޝRzW&=;J������� F�b���tL�0���M�=S� ��ؽߌ�q�X ��PVò�� ����b'ulgdb��H+,L��#�qo[u���B�	������\Kj��-�ΐ'B-8!FLBJ�nl�tq�]�pIS��fQ��]���V���S3�����o�vP��
<��l���R�|$��D<b��GS�N�'�*��"4ҵ�)�Re��+���@�s�q�L����YXۺ�ʹj�*~������ �'Գ����z	���Beρ�`�T uLE�����v�Y]IBİ�	�YN*(6'Ud)�����+L	0} ������Ʀ&�4y�S"k��7���`��,q��啕��-�F�P�9��$@���0�W��sn.Ĕ�"@������eiL��{�T�>��Ō��=Ý��Լ�9헔��/�r�D�d9��V�M�f�S����у�%��Tj�O4�M���K�t0�?X̪����y�T|5t�O�	w��eX܅�!tPYa�o�����x�ۗO��9g�����v���ꈣE�@j�s\~�E{��(B���q���+)]Ո��ik��RQ ��NԜ�ooF��(�75�8O|��1bfH/�,������|�������<��xa�Y���ږ���.�J�}�x��%���na�!���S+舓�'��4��	ix;����!x�0�c�͟�JʈC2��ڿ����X;�G�������pq�d�z�EIHH�Z{�1 �eR�r���5�Fv�B��t6#+)�U��ٗ��y˖��8�p��ͱ�7H����}���G��� o�p^��(#m�V��{�6���?A�]�狘�� �C��N:���u�������s�Φg�|j̕z�@���uLQ�?4Ѫw��7f	�ׇ��B�>� ��[þ+��颬�r_����J���V|��0!����9�v��Q��@� Ć�?ӓ�N������Ăl�^{_�oV�N��|Q"=%���`2 ��
⚳�]8��Ha�vdK|���=`I�������"ζ�QW .zE�L�{1fp�ܼq�.'�@�:J��OPZ�4S�p+��]pPG.  Pjy��Gk~���#c�&�r�4$9�º���*S��`a�`�i3��m�9~�(����v��e�ܿ^o� �����WRx+dy\� CQ	�kQlı�İQ_?�� �){����r\?c<�RL<n^'�F������Jǔ�yC`��qdR֍#��L�*��Ȥ��hl�jK�f5	�`%Lu�A8p=�5`_�c�����՟đk�$3��mB&��1�����D�=�-ٺo���6�q�TKQ��B笁��Of�u�m�:��R��Z_�=�\��R�Z~o<�M�zzzȜ���tX��3�^���7).O��.�z�^��:��7�L�,^����λ�ǁ�k�T1�9��t#�i��Y���9�M�C .�h+��w�@��R�b}����/]�$̴`�?�v/ƽ~��<�r"S����)P�_nz6T9�l˔���)�Q�O�j5V��1o�?�CO	���Z��m�4c(VT��1�=�� ��X��c��lͽ�ɨ/�
ث[-_����B��:��+s�j5K�@0�c����v�7����U}����@$%��>�2�a���{��o�������(~w?H��u�c�4m@����9o+��ʖO��%q�_����-'/l����[I�R�V��Op���46���l�-�v�gD��}�@�"�U�s(�]�߰P!�T�ܳ2����Y���dG���F�Cƚ֭'^߳IF�Z�n��ߙۓ����C��p����X��FV=3�� Ny~}c@�8�8w9��*��JG�2��c��nDM��[�l{���g8��#A��<�h0�-�G�,b����nĀ��Λh!�D4�*N����j��	�����,
�"��i�1��$!PRۖѶZO�W@!��~jk�`�s�/y|����92XP�Ķr.�����{����S��������q2��dOc���O^����T��˺A��5��g+I4j��7Dm��Kũ�>�V�>n��ʙ� ��J��9�۟�?��l��' xu�0�a���|�a'T6�	t�r���5��Y�dh�
u��U�2� �U �Lx�A���܃̅Io�s/e�����)`����5�q��o`psO��@+%�"�f�O�i�؏o�n	O��X���1�:`8�>JP�!�('��/�53���yl�/U��t�gg[�+�uNS5��ˡ�t�"�~o��OgzD���d"n�P;E�B~��؉�,jݞ;U8[���@��LF���u&�W�8�gI���7#�z�⓬�ڗE�k��]>J�%�*���C����N���	Έ7���8k�sǝ�.�?�	��u��=�*�:�)���sz�Sʿ��v���-�D����4�̈́�Ѻ���#0I�`��F��`X��.�w�7U3�|#������I�i5�yb�ߘ�o(c��>j�H\>�������|��P	�Q�>�#��-U�����~��Eҳh� kDD�NT2T���7C��G��/��p��<��������Н���wDa�K!�$9J���b*���ig��L�/��N&2�9K9un�]����O��!�����W��E-���-�ݭB��"�x+�2��#֯��ך��?`�����!�gc�T�l2������Ӈ�6'�<�̓\>˰r_�]N�E����mnh���ַ�R*�Z�dxg�nrw=/�4�~~�c,`<i����"Y ������e������n���o�.W�I�|X�:�(��/N�)=�L���+�*�����R����S9�I�ڱ[�,a���W���Ŝ��ڳv����������t����Q�� uÄ?ҕu�����dr����¿8��X��r>�Bb�ܿ�"֘��g���Sfv��g��%�u�h�e�VSH+�]g0�'QN<{���P2�{!]\k�p[���}q���D˸�o��[�C @`n2�p�Z�`v��/¿m0�ܿ�ȭ�E�o�����{�xF���� ���6��u�j����eF� s#�T��j�EY�G6O(�%���p٤�;fy�YDIY�	�ͮ�\�,B� ."��'ڈA���gj�w�"R1��mf:�୪�=d5����u\C��&�nDC��G��ܷ7�6a5���<c���	���o�s����R��T�gAg�ao�h����n��RR7�b������`�<'C�����,eZ�f{Z&k4��ƛ���{��w��%a~Z[���g�m�I��#�UƟȍ��&MO�?��3�o)+q����'����G���_حq)�.#��'ড়؉A��ِ\���'�A����1�����[G��f �?O�6��ۍao�K�t�q75�X�N�mY{J��W����*+��x��?�מX�)Y����6&�$��[�S��s����8���A_��4m��qd0N{��|O�� `^�����^H�~��Ǉ�Őܹpy>W��Të�rw{�7qh0��V�*,:0�WY�"����pЈic;{��zV�c4�*��C�B�Oا���۵�|��7�8]>�!�
:�yى�!U.�[�wr�'�U�L��\r�kL�ڸ��R�����qn���n������B�ۙ���/��۔�g���A��쮷�k�G*��e3d�ʫ���d��,��}}DP�p4e#�ݧ�蔂��r��YF�i|�:����
Vm�]?~�!��yh��9���~��Ή�	�P����2�򽔏�:&4�2�$���t����B#�t����$��g]�p*��Ơ����J��ɲ%zJLL�O0����v0;pe���a�mׅ����)��X"Av��U�/3�Q���̪�Dy�|��;%*)��ˆDO�qwԭ�Pc��[�M���,,���������� �g�'T����T�F�x ;���)���P^����ę+�9a
c��)"���@i~{ic\�8���U�j5���g�m�F���7�o)��*�+�[�:��Dmp�<oz�|(���wf��#SAkAi��ot�<q���6D��4��q�#��y�iz��b�o���'�Ok��T�RL[���kA瀕��Pp.�$��P3y��>ѷ4��ҡ%b��¢7G�*���r�2��Gΐ�!n��tY�8>� �f4S��L�<�@��t�"7�p9b\�4`�����q����}��D��O�.gԪ��l���!uL ��w��N�C�^��K�z/��-���D�k"%S�J��*��toٮ���c�Ϯ/��n[���*�.��~��=�C3MB�"Md1���Q�tS�����u'1L�#���Ƴ�_�=f�h���@�h�'�D�0�R��ܷeOG�֨j8�j�5�V�Oh��]:g��[��+�nZ�Tc*�sՕ�O�D:���3�H�7�|�Af�ҩ�g���`��u]����*bm���%qѶS�ZW����`mf�i�[�W��zGc��6K��ۿ[��b'��3�%m���w����z���S�E}�:LL�)��x2��Q��Mao��(}��p�nE�!��1�6wҊ:�{�#�5=�eS���$M�&�/�7:p��샘�1�l��N����%�����մ8�.?�ڐK���Yos3&=60��9v�!p�}����c��
}���<�5#B��K7�X�k�e�X�^���Nl�n�ȗ�����ӄ�U��NWJ�/�?(|c�: ��q:NxӲ6zR��>9��Y�'Unj0�I��uF3W�WK��?�wi��(w	:]WjZ�}lb!l���:*U�#�j�
05,���
vz�=��јK� ��h�X����B��,5�il����4�#�?j�6�������{P	Pm
�
�.-ݙz��ȍ�Ȃ+{��oA�u);*�BDk��x>:��2g֞�����f�$�:���}q�L�0q�])�9�g(���bB(�X;}�u1�ˌ�Se#���Z��/J���,+�Ə�].zf�T>ݰ#)'݈;`"�V�Q�-a��B��7���˪<͢-�2)	q��+�'�6� �5���m81��A���׼����~b��_/���`�z�+���ׁ��yt:�R�/�b��Ǘ"���˯qj�j�Xr�v�m�WE��������cF��	�0[ݥqt2�a'���m/g�u߳�Y/�n`p \�$h�c�ӵ?�&��>����]*ӤP�ǻYs�q���w0�mS�X��y2)32����V���y>C�҈���(#��v�����=��B�o��_�;�&��vYS�C�J�Ȧk����0d���$��$X0U֯Y�ۙ�-Z��ft�f3���sk��W���H��vMx�9jFqch��;��� �����׈�����,�\�^qQo���Ki�3b�I�'१��5�{;�Ð���]�ky����F���6Ow!I>����8+�3��0��>Q�>
A�RB`'\���)�%�П��j�7]iX�(�x2�	΅�ZX�.q�И_�wa$�Ӊ��m�M�|3�����S	���F�;9<IXDpG]y?ɹ���ڿ���q�����7]я�������|�7v�bDŝ��4�B�z���g_K�B̕���8�N���'6	�b��Ë�2��1R�o��KwΒB2SQ>jE��Z��<j�0�D��!��&IIc�:�e�i�9B�S6�(/�Ǌ�݊�+&Yə
���YC��0���W'����p(�#w��Z�W��7Xx�t��w��w�����u���"�?�n'gկB��UHi�T�������T5���}�[�Ŗ��po�\6\t��@�+�̩���L�渡� }�cEq���(�kK�t$���υ��� �)#lnT�e��7�T�dl�5�#����l橫��� ��A��uq6Qe�N�
t(���=3��r��=��i�s�%T:s����m��*uף��dl�����1�Wi*��	������n��>�s��5��@+jGLL�Ȭ:t>��G �G�u�H��H��ǥ*J{��ns�9g_uciX�1�����|á��~��x�&�p�F��@�q#�Q�3������-ш�����/�*�Lu���a����r� �(�Kj};0�'�J�fd�O��pb�qm2��ni@�^�ؗP��+A��m�s�j���2�5�	]�|8�`���l.�����������eF������DⅮm?'w?��[6��-����\�a�^Uj�,t�p"PP���hr����x��8S7�v�#=/��Q�p8iTu����Q�8=ϱ�w>���[�#LsW���X��D�
Ê���FARH����Ȩʢv�N��ΰ	�8x0��L;�Y����������b(���g���4~�;� :1}���`aU>˽�ǎ����/[aY��>]~U��ok��6'�<�<).�����}�T�@lv��l�����\)�;{"A����CA�À[_H�������H�UM�f5"�Z�h"�>1�0��`5@�����e��"���w�B��� ��V��*�c��|�!�Mq��[�ݿ��w����5��v�:�yA������$�OZ���
�T8����EL��f��Wg��(#���J&P\9.o�k=�˩�v$_�a����]!5*)��9��A��v���ee�ƍ�V�eW��7�cw�5�ml� � ~olΏ ��k�̢+�8�'�)n��7>d���A�0��`�&�s�X
r��8>n�6�l����e9s=��,�b~��xf�'�wk�.�|f-Z+�g�fΩˣ�-�(�O-�'��+�z����Ƣ��}*T��/=�8��K8�V����q�4?T]�8�Ɉ2�A�3�,7�_����+U��ݹ���g�y545A��6�ʥ=��-�h��EMC>���ul?��ѓ�yI�q��D���X��qF��p�%����H!�Kxy]1����h��BF���I�l$|FE��u�:�Wϧ�1���s]�9�vUt�:���
?Ek].��%zk`��_�`�t�����*���#���E����s��A
�JZ�n��4�@r���ܠ��E:5�թyyG��a?�?��l��7�[&��bB,;-D��䈶�>pF��JgR녌���؏��]"�.��&�kV��M�Iz-o�&.GRt��.�����B'PCb!��(V#��r�x	o�B	w�y �E[·&���`@@�:����)���8U��t���c�~1���R\�x�۳�O�`�&J�KH�D]=,��(UJ]<�4_�M��:����v����^�wǑ(�'��n4G*�l7�U�+���>	�ȡ�A�]9Jj����,F����,;�i8�0�⁇$I�^�tuK;:H����X�6l���n��ެ;�(j\��G]�ZYO�a���m\_�<#J#�d�EP�x!�]��/d���u�s%����f�6^(h��!g$DU?��-+N��9��H$U�ʴb)#�BA�e?dZ9��흡tĩnEE��S�����(q���1��	%���PV
&�Ut��qO`���]��|#�e���c��VYVOA������]W��W	Q���\�,�9��b���ѷ�Ñ��[�7!�zbz������on�|��#S�rYYL� %$��&C�U�͎�?$����m��1����3�2���K�"�w���}��$� �DF��b(L�$�I}�	h66i$oU�ܸ^�1�2�b�C,Ku��f'ֲ�k1�4rR��C��28v"A�ə_,�r-5�%�f�����v�뢸����*!V�Ck�ŗ��=�Ӣ���ց���O�Qy+���2"ϱ:c*r,�<M$k/�6G��G�4�E[�>���'�y ��C��m��f�	��o��{�EtX�Gp�Vxb���v#�j�A3��Q`��)3F��r�PW��%��`����W��YN:����cT��B2Փ�?���3d-3�f����5�[t��w��d���\�,h�:8��ao9�� �4�nEcC{�Ė��PGo��wt��tn��(��R���c�*��y{~̱-R�*��!�r�-l�K���w8�;n{c���dX�Ġ���U�l�kQ�G�D�qxk�2�}�Bÿ|���������HY�,�G$P�"..����k�H���$�2���P��K���O	�\������]N�[,��z�/<���	�Ykz�щ�n��&;�2����.��ǖ*�an��X��,���u5���d�4&@�w*Ǒ������p2�����Y៲����T�v
��BF���킖-��˲3��^�v�}k~�X9�����ǰ4���m4����"2a����e���@���9����\�t4J��0�Ԧl��S���-��ʮ|l���
>�3(1SNgl�Ȕ8q�i�D���6t���ć��EuO��'�^�Q�Ih�}}zOe!|S:��2�*P��P;%������Q���,o܀����+0ff�% ��k'S����}��Ӛ1����=�ȕ��oN�����@����N)��v��a��~.�Tl�Wzk@'66��I�f�u]~J�򤁃��U4��Q�� �J����R:ā�\G��9���d���dg��5s])
;������W���7P����J���^g��B,�G��_��)�쏼�ߚ���B�O	�9�Vv�v|x>]	�ė�{�tXy��um��w�;
ل޺A&��M������|�Z6�Tx"x;lb����^�fh E��U��8fl'\��`	�����V	�9���'v�˝ ��{�/�l�?a� ����e�>ʒv�c��ł������%Ý������������3K/F3Vy��m+/�Ba����w`�O�c6LrV?~�( ���5q�PY�յp�JQ;��jc�/�[�)@ͧ=T9`�ݣZS�\��j��R]�(��,�%��AxY���%���_jjԍ�1�)1eee-��Ī�'��C�W�v#�8�-��OR��;�a3vJp0)zS=*�񫯭E���C�#����٢��mC-I��;�_[���g��m-�-�q����S |ϰ]1���-+�[�$��39>nj�0[n���E��FF��˭�,ǅ�v���I�3�[��ki��y�ѡ�o޲�&:��=d/��?)�h����kɰ-���:V5�Dl�?2�m�<�2Q�R�&_���E���y��ΐ�85#�����a���~	�|C]�ko�s���6r�_j����}K҈d��2��eu���'g�B:ǉ���v���)�z��A�=�����4(5''���S�����_lRc�L����C��+� 2B�����e�Bג����y��sl�&pq.�=�xSS��SZ�8@|���q>B��WtNɩ_�6��o:�S��� �q��l�^0��v��W֌�ع�=��i�r����u�����?��U������`�9��4$Xh��*k.��u|W x���zp�{9�j��E#gM"7Ƹ=�a�2E%C�I1׮Mz)�T��	�N$���ҷ��m�4��9;�3�)�s�%�K�����1�+#��_o�M<wBNhh��P����T||�#�9�6�e0�>\�u�&�>�\��	��.��i���rv:�������qX�A�6v�¯���/w`�w*a�����e�����7o��Z1���\&WA72
���;r/��~�>3��-�F�!�Jc}�S���LQ��m�=�/���7��4�/��*�4�5 ��Y��4�����;馿E	#�&l�,��C:�!���FN}9��H���

ʇjuS�6��f�I9%!Զ	Ѝ�,�_h���0cQ?�K96����!��@,�!k�#�S8�:�(݄�����Q�&ɺ�+.?t�d�ϣ�d�_�q���ظ�����U�@8��%!�[�Z5,��gyH��<7P[bk���{$o����I�Ǌ���[�!�}�!��:p�ߔH�0	e�{p\��c<��8�:!����,�k��P �OxM�FE7j��y��t'����kPw�WĿ��>F"F��1B�J��E���ǿP�J���FP3�<��������˧�n3+�#�ɀ�an%��˲E.��iú�j����ţd��F6�#E��9a�_����8U�-Po�:��)mG���Q�.}'쭫�J�o�~L�6�@���ύZ�q��.C=���ea��?���������[[�37x��hi;9��	yy5Y�Z��Ӯ�F��G���F3��~�{;T����.ѫ s�
� R=p�M���az�e�x�����s<�/��y�� �P��[�J.'�j<H#H@���;գ�4~���T��Q�ttt�����"[��oHIъ'_�`޾)���=	ƁN�O�X�A�.��2�� �����ǯ��`Oz��ս���v}o'0�|��˟	Vfݺ������{%A�x}���>jUҠ"P�<q�^X��H�'��7b�%z�b�(����i��}{�OO�W�$����w����kr{6���N&pqC�*M�60��:�%�my��o8�Xh�Ā:5��dK���b��
Fu*� I�&���K�͗�;�/Q�%U�ᅴ�'R0/��D�!��Gm{4�8�L����>�V%iѣ9b�Q�	�A ���a[�SKY���=��I�)�����ܗ�̰@��Î}�6���M@�Gl��
v����yf����"��uЗm���[	���z� �/�7O���HBW�6�V�C2�x�1&ia��9wR��k>�A7��ħ��"6269y�ݝo�c�Bk��k*�@��+�$����*3��=��.+���D*AB@���i�É����N��}���� �p
wEݓ� �4���"ͥk�lA۴����1K��Z���'"�d[���ӰI��L�4���Us�����W/ը�$���OG��>*�HO�=+2���b9�U��go�F\��/þ����U�f��,P�i�moo���9c������E��������o���V��9�Ov���(yY�Ʀ�ϋ���������?�}Ǌ�s��s����0����$<�m�I��H9}�(�w���,��g.�)x�Tf��)����H�f���奋Z��A.hF��b)�(z!�S�i����P��_Mfe�J=x��rD�'3N�۷o�߿���|>�?;>>v�8���q��e2n���U[^�q����ǰ�-(#�Y���B�V�����8Cj}��3�x�p�">̡K=f�����o�F��ǔE����h/�>`_ߕh���=�^H�����]�[΅Ɇ�]Sy�s����P!�22>�0�h��p��)�h��4�� ���O�0>��*��֕g���g���]@��X���_�,B��U��w+�{wcE-n�<����N�m)ڬR�@x[�\�` ,hj&&@!���L�-��iD8��R7E�!t���]+��2��$�A�w��E�:61�(R�ӆ��R�1�.R?6���18r��H%�3��g,�ݏydF-���T/D�{�<u���ʦ�I�M�@�����y�t�B��	k\=��n�%�т-u$jc! �Lei�*p��XF�8�g����xx�S��"��>�Wh����-n���8JZ��H��$�UuuH�t��.~u�Mmc[��|�V��h�c�x�������F4ް<;���]3b0D�f<�>���W8�j�����)fX���2�"8)�P�HI>�_d��'	?6�yӌ�X�<�K�����G����q]<��ߧ���1l:�x��/�A�,X�7����T�;6�ɲO���%� 4�!A;G�W_�z'�b)�����-���N^�P�]A�"��;K�ٵR�˵\��)�7��
�i�K�{X�#�t85�v��W1H����U���"�M�����~f�0c��R}��C|��#5���AǓ�O�o�l�?>HR���	�l������Ô@b� ��
��ELqH&�ݰA Dy�[���@�?�N�l٨�=������M\:��F��;�X�'j!�XU���m�pQ2��#��%M���?���.(Q�<\�EVAº �>�Q���&����#׏�j琊�W&M�hy|���� �N,��c��S�p���m۠�&�C	Hܓ�C�Y>ĘK�Fm����)ԛ�Y����w��Ox�+���b��xz�^6�'L�YJ��z�8�D��ɑ���8�\!r)���1�.�(�s#�������-[�B�|���fξ.�G��MII�H��olB������y����TXV�!F�p�ԫ<s`)w�1[lv�D&�����G��B#�b�� Ɛ��W*�!R/n��Go�~�sE4�T��x����X�!��s�k��UZ_N,ǭ���� 
}jv�f.^�����O�/?�S���vD.�c���C��%���_��Ἄ���%��n��{E:�w�Z_�A(�E�#�q<�{oq(�	Ĥ�R^*��`c}h�����8��+0.;��nmn:M�`�f������>�J��5�_ȶ� (�E������Go���}���F�#����EL��$�G���*#������!觑Ў$��9a_����lq�X$#L��1�[�:t���k�Ep�A�444|S������Y�]��}��gP"��g$6�&n�2'�dR�kl�^p�1�X�<�� �IH�0����ǀ��a?M�#q/<1�h���J��h�]��۟g�oc�5���̀Q��<EG(g͛�G�A,WQ")¿]7�k=���D"��u8���Wﺺ$p=vG�N�U��v�-��Q4��z�SI�L�>�hW���Z�>g<F���:9�.�h���l�L�L'qUҀ�!@	���}���p j���ӎ�?�i=\���	�!����\H��oe�+�*��H(�(����R�b~��t�d*ФbW\>¯* o�E�>t�$%�P�(���+����Y�-ەh�T8zE�����J��o����{����E�M
�P��3?�ΉX�\7�*��!K�6Qz�RZ��d.G�K9�u���֗��_��ͱ		�?n�?4\T��^�C:���[D��F�s�n))����)醥�k�o���9;�f��ĽwƓG�zRl��}B�r��5}2��9�=�j
�2���"�����v�E��E2�^�
r���\\��2�C���mF�ͳ��j��m�Tw0KU��s�Ն�n	t8aӫ��xY����ÔSnbs����kg���#$�����)� �r����^K[����n[j��������sI@V*�XX@�G-'�J	�.�
�I��c���a+����)w�%6��*��˕r�5�޲�-q�3�k�G�x�?��5Y�1f��1���z����`B���ժm�.�6A��l��B��=������RRR  �ZRX�a����.t~�j�zbp�BT��	���k��{���3������|x=�3�a��gô���!XV�	��1���k5f>�[�6B\�JToX6.����	H������1�u)�@k�p.q�I>j���������-|�����9��;�4v]&/�q/"�ͥ��1#o������B��\l�$�D����N�/�l�������8tj��&'+Y�1�״xh/;))� ���e���!#V�n�mR�o�S�ʰN��Л����#��*v$Z�i��MѰ	9��
��QQUF>�O����̚jj�!���X���\NP��'��[8���q*�Zen	b�~�A-2}_�z�+�%���`�g�Y���|ˬ��u5+O;�����w�Mu1�����	m��߂F_�t�?���sx�^���[A�al�#Ҽۆ�N?A��/���(��'-ԛnB����>~� ���d�Os�� "qX˨m��o���Lysj�?,�
z�ʕ~���.|��;���Z������x��7��&n��7��S�� �`�&�f⑹�U���)�ʧ���<� )}D"�i��p>����j���p��ܔpc �,<p�ѽ,�VY�d��rn�z�L+ ��t�i�0d_YCAV;��Pb���+my��Ii���h���G�1�Y��u!h(��a��tϵ���@�'���� ։r8׍�넞]�4"b�
]7"�+v� ��!wܰBK�T�>u�ݖ(y�������A���3S�|�e��6�0.\VB-s~����G�l$,fZ�/�#XK��m���M���$��/����N���d<w�5�x��P��%���v��X��7>)#c)#�tb!��Ce�Б�8�����d#��8 h�v��7����)$߽9�zӳ��ړm�7�&��h1�I��|w��}��'��A��{��cͿo����c�F��:���M�b9�[C>v&�/�i�5YҀ��U���Æܗ��=^Vf�{��qwO@\�����ZE��\:xp@�t?�^�����d�W��x��B?G�}/��]Gk:�d͹��v�Xg����iE^�R�0������ąeۺ�鰳�KC8�%����"3k���U��;+�	��c�H�'���<��'*�)�d�v����3�A��V�R��@�xA�+f�ԙ��P߼�h�}m?�N�%�?&d��)�]B���Z��l����_]�O1����A~��4O(^_1ükP�=�	��1�ñZ�߉��;u�5ݾ����Q����~WIz��h	�l�5F�u$�����zɺ�#��Z��ʼ������h�T��&z�M}O�:΍��q��7�\ߧ�S�K�IYJ��}A-�!8xgUW��J<���zd
#��$�D\��b�1�k\�	��&��S��8.��Z�wm��й�$�&xlɻ�* ���1��t�ngVv�]c��q�)�t>�]��1f,��C�yjh
���FhjV���}�Api_�.	�K]�����"�3�ӊ���0����&������?���R����|�fmHL�]�-�o��_�[��jm���i�U���e���{����h� �lnN��U~�)�wL���9����вr�8�'%؍u���SsHi�w�{�:��i�÷|�t�������$.:�9�ׁ��w��qv�=�Q���j������˲;D["X+V}�>���iP���iP�W:1މ*@2X��K���A�ȥFp�?��9y�L
������o�����aGmm��c[�7c�x�*�SN�"��a�w��#%�U�Am��K� �u���]�>/?R{/NnG�֛D�!mI�o���}Y�i��CvK�Z^��#s�7@9=8N?���z Q6�RY��F�2���(�7\�7D�6�)������Xꡏ���R7-��]���F[�,������xh�2k���Ӆ�b���[��%��ʅ.!y�]z`���Դ�k��Ca�1���lD���p��LΑj����X��Ǫ���GH2v5�¨�K����ӝ��d�Т��Yk�Ē���F��ً�w~�8��=����%Q��+O��;������/��؎w��A��E��XnK��f�`>ͼ���맧�k/S��c���FET�^	M�*�놟A�˶F�-Qg��g�q����ɢ�?�q�M�J�?�(����<ؿ�
[�o�R$66��͘h��0Tz��[x���	�Oɳ/I��^�'u��������ZQ=�}A\ �+`�l�/��4�s6���8��=��O����J좺�7Z�7��O�D��2��������*bg�s�ta7�CA�`����@�*N�d�D����I�}�ӵ�^�ˏw��b�Zk�mH��'�yF��7�5ɏ�}��
&"���ʎ�V�> �=��uB,Y:R��I�����>[��Y=)��o���g��.�UT��:��w����Q���?�0���,�_��wO�/gz�-�]�g8�`_�qyz�Fm+��?JB;���������:-��e������N��R��؎��,�T�5�;#Q�Ѫ3<n���M����WLV�u'�^�"� לiJ�����{�8�p��ewo KQ��ĮU���f	��8՚����ۅ�K��o/����"�$�D��a���>�G3��u�I����)HS�ʶ���#7RR6��粱��}���ɷDCb�dz�j��Î����x놠�>�_��`.�t�tt"��8��\S������L����|{u�2�Nv�ۤ�s��8u>�tM�®�h�څ�&��v�$|*��ق6>���×m�_�*-�1��c{���"��{�l;NRh<�C�)k��v,���eTu��z��ME>T��/l��M�@}�J�%��+.=폯���y��bM�f!��S�9?;��W��;f�r@:���Y9ġ��9V�0�0])��c$
����U�6pqnq:NQه_�E�q�&~s}K?����@���C �(�p`	c2�U��,�`�ɥ����n
�\8<�S�1;���U�����K��3A�l�� �2�K��c���g���kI��,&��.(T�$�L(����6��������ʄ�����b��ו�P��C��}H��[�����2���=VEp ���0^�	��У`w�C�2���41��7�����#^��������g L�:��U=��yK���G\�ܦ��H��i�`����-H�2�>5� E��8h�p�E��%���scN�C�"�Pe$A�g�&.�HI�맩x�L��؆��)�YyU�(bq��W�?�5��M�R,��"&�@��	;�1��m�8.�4�%Ng�K��Ԃ�y?�K�RR�w���1��mO� +ϓ�
rH��:6��r�a�Ɏ�	�Kd	?s��.��̶ʞ�9�U�;D���=���ȓ��)&�G)#$�G�	��'a�� ��Y�R�zGF�������i���׆�/Y��+rJ�����w�[q��oy�?J]����u�J{o���P�0,���8�i�m���UJ(��G�T�0(�e�u�ቻX]��;\�8�I��xS�q�����p*�Gb/p�x�&�!�b��<O��kA:*n>9f9Rfp����ɰ[�X
�y�<�B�a�	�$l��C���f*���Q6B��4ǲa�ἁPV���6�i�ǆ������r-�x�ڮ�.�˫�cǅ<��vc�a/]�^iJ���(���	۳������ܼ�Q�	���`��t#��&���Jk��P���MVD0h���8�E�C�n�\��5_s}�s`��t&��@�cg���E6����>��Y��	,�0�>���t��ڋ��-1x����¬p�[��l��и����P���5c[��6�.TVW���Ǭ`��X���� %�^�t�Ͳ7s���(jL��}�u55�6:��ɜi̢�a�ftM��f]k��gAH�� v_v7{X@xl)�����s�����*!�W�+�(�ڃ�!�!iy���l����C�RK�d��k����!��ht��+꺇�t��$����m���[8e�S�E��`g�+LV֮�?�c�Ç	��,Ë́�O���r���D$��+���ß�z�� B����0��<Kq7pG$�I}�z|�Kt�OYW拉�����ԵC=1ya�!q�~��QX1��S���Z0�!8J
Z5\:vke�D�����=��a�PR��A�TZQ�	2G�`o�̯_DA���`�S��\�!���uP�Kr8 �=ѽXm�L;Pvt�5�io	��P�V1��%E&�q����wP=
<L��oF\��g��?d$�`�E1�q�����P3�s�ۘ@!��R�u�&���T�Z�MH&���s.�Vu޺^���hgFM� �G2K�F�������}?�RY�N-!W����+���ߐl���>��=]����c=������AtY�U����ESo� U�O�"�����>�M��~FK�e��+'ȕz�Vg��U�l��g*��ʈ�z�#�������1/�������=G�N�G�Ig�`��b���:'W�n���QM��T��z��|��o��bcWUUv?�
P8������L�<26�r�f�7��~Ch�s��Y���|��B��C�f�*>�ojK�7|�_QK��|������>���8�����{C�ׯ��d�sO���q��U�5��a�;������>�R+�_��"��K�x�_�i�e��9�_����: <���ֹY1)�Y�ѻ��DM[�����>�o�3da��81sǔFn����{�[V?�I���/�TD���`RP�ny�v�B�G��h�FV��^��Fv�Tk�uX����h����S�UVĜ[E��r\��ǲ��@�0��dAo)�JA.
�d�T8 ��i��8"�˔����r1jR�]���ǂgO�����ӏ���OO�\Ÿ�C�G�6G�6c,NaCa�ø���a��^��﾿hս�,��t($ddT��Ǳ�e�W�)~,]�y��k����pƚwf��]�>�8��~���=^�d_�ZX��~u�Hɗg��p?:r�08%x�grk��V�3L]��$8!�i� :x����~�+����d���[$S{4ɤB.F_1#���VR@�����t)!>P!x���~�F^drv;�QQ�Wxֺ)f���\��Ta#}Ga�M��_��O_��{l��.�4�x8�|x^yO�8������o䩻]S��z?")F�I2�oe���cyT�ЯUh��M�76!.mJD��
\��� L)�[/�TP���S@�#�����"�"z��C?
��V	��(S���_�z~�"?�ˠ{��d7IIH��_[��(�2:p�����#5�P HII��qar�����*�sw�	fcȋ	�H�j�N43�D�g��>]��M�y�2���l}qk�.П�8��v�i-�* Q��h����'�X`�[�]K���R�p�V�!`¶��&v���0�I��b�+6�_%BA��q,^�ǢSLߜ��Ǘ��Ă��a��X�
�����.pr®�UǕJ�X5a�*��ke�!���2@�.#����DZtyi Ke.} ��2�R��}�t,,ż���m��{$K��I�L4�K2a��|-�IB}"ą�H����Ni/��eUUD�S̞T�N��S��u�B{�i'�R}������>RO�+�\R�򒖗\�G�7��D ��k�����`
��x��Ui��`�~y`O*�+S9%q!>����ё���q�O�c��vŘ�sv�ՌS���T�1A��`�a�_Cs?V�ck�$�V #���l�yn��~O��+}�4Z� ���O<��I��a=+�+;��I�u��ЈD�n0��F[��U��8gvv�K*7 �!��uv�����U�I~8q�ڌP��.U'DZ��N�BtL �^�@n.��6O�N�x J�S[�U�{�;�ϩЋ@]���d�j�.��)[CL��[�PE;~�(�fj���<՚Z�WJ����>���p	{�+��n��Ԋm0�=������I׿#��2�j��A�G��V��8"o )-y _y�Gx��O��m���qb�V�L�7uie�Q�u|R_m�#����d�.��7�Z�"��Z�̈�z�j<�����"��ñ���k-��l>��s	�e�Jn�QcN������_�k>�S�ο����å�Y����H� �|t��j�oF8�Z�r`����􂧷b �L�ʖ=��)�#�n>x	��}GMt�wʬ��P� 6��e����K��� S#5����ZקnA]lX�![���7�p�~O7f��O��;���X���+7b('FX7�E��������^�����,x#��2�d#���#�Ev�m�xT"H_�4�4�8�ݽv]Yp��.b����������)�\s'}���m��u6�������5k��B�p��)f��F~����}u�����O���pϜ��o�Vz�冭�M��|zFgO��d��%$���]�����񛮚~�t���0A"�P:�Xt�o��y��'��?{�64��<�����(HB��`J�		��ۨ^��M��k�~��x��lN�_"k�F�xD�$fm�g�Ȭ�4l+����16�ga�y}�#��	�uMR$�Y�=��Qc	�-��pr�����;5n���
��� [l��_e�~N�=�X�Q�CB�FVY{���sە_W��!�Ƴl��]E�2?\`����f���rʰ� ��w�}B󃼨�|�Oΰd�����f�Ɇ�-ו8�e8�|�K>��{��R���c�Zu�L�s�Ȥ�����GX���~��_��o[\ɸsy�^�h;7l�T�g���Y���%���fW;΋� e0����g��`���y���>��p	�ٍ�Z0�KwZ�z7$�FwB?�:on28ނT�Nv�h���#��;7�sZ^���6Ή��p9�;B4cKzצ�)�]�O�&i�?��?gL�-�@�٥S������A�ROez��c�o���
�0qȀq�E��e�`�(;s��g�@���'#Q;QrwmÑ)�%����� ;�ܾ������`vd��AB�_6�h������1�6'���z���:-W��)�j��v�_<�FF��b�[:�?����<�Ո̵���[����~~+�O�%���lP"EY�-�7�O�>d�.�s婢?j1lkw�561ښx._b�U�4fڒ&!����`?R�]��r�nȫ�O��~3A�0/�DF���j�N�T %(\t<x��9��?�F�nJ�T�SQc��؜��;���.�f43G�����,��[�~���I���R?�o&�f��,������G��F�f[X� ��,uoZ�Q�63{��O�l��FV�jR���F7LAy�S��o���((���G�-����B�N�	�D��x՘˅MR���is��-F��bXT�Q u{�W�6���
ϓ��L�:��>t��o��E�ښ��÷�����yhu�O؎N�W��ʽ{�T2��rP���Z�r����v���8����e��r:�0�1>�������X$.(����A� ���@��Ը�3�Z�ؤ��!Ez��86 W$�0,�ώռ���Ou��-"��Vy ~�	�K��ű3{c+�I�g��~s��x�"��9iK��v)�yK+��@B�@�C��y��?ּ�(�b���To�s	y����ᱰJ�+�б���Qô(��>x�� ���;�X���'�L���њ�jGޢ_��H5��$ëQ�O�.��h���e��-<q��w� M~��O���:36�v�);*��77��b���
<������2��a�ʜ��b"��JF"���,�x9��w̕%	�����hݱ魖	�C0Vi"LVA
b/`���x�������P��S}�Y~ϝ )�R�?�F��@�t��"�P9ҫ��a������Q���D�6�+}j���1���>��>!]���m�뢂�+��]�yK�e޾���.��
�,��ac����WT�?mz[��O#�*�[Ⱥ�P.aн�L����_$�t�3L�#�$���W2��H�xOWEr��v��:��U��\�s�AdVS� �ߟX�}Ԗ E9EYQ�#VL��F!�uv�D8L+�r������nhT���S��W��(W��t�t"o���<p ��L$����LNC�HsQ�wR���ԣ�)U����VJ����1�6u�p�@���&^��Q�?�rD@*?�ۥW�u�M��;!K�Ӓ��%����m�ԦX{�ɐ�y��H6�_���s��)�a�A�d��=�HMi�2��� W�qU�_% ��;�R�{MP�C��67����wg��� *�h50R�Z���*Ȏ��\���er1Ǎ7W�e4&�O}Œn�w�x竏�lg��crv9S��eP4ꂭ�w������WM��FR��ѝ��&Z!v+�GwH.�Ų�E��X����Z(�ӥ8sbߗj�f�(�3U���b�K��]r�����;Tj-Wּ%.�Y��0�曜�'�Iٵ�6����Cf�x�8k�����8�*������ ���PC��3���,��P�s�ꆌ0G�5q�uK�{_?4u<E%��c����raT��I|���'�N�\�'�ް| �:��y�y�~э�����J��/y�{OFE��KP��&jp��K�ʹ~M�3�nB�Y5H	�Oi��6�U��|�)���\�5�<�32�>�G��p��æ����RKV�S�q�R^8<]Ykm�{�YkK����=	�����<�V1UXlާ�}?�����#�d��l��g����P�����R��q��U�
����f�,��V�d%��^s��3��� ��,�V�J� Ù�����7��=���L;��)v��6��(�ͬ�&D�N���E�F��������2d"WքH��o�=+��`2�����f�(�����^(K�G��0)�Y������	�Et�W���Q������n���wU�M�dٳ���-*��D���IOqӻ
;��K��:t�<��^8��l���~�� ���?j�4�g�
�|����g�� ���c�2��ek?\;E"V�́	�����-.��W�c��ԚU#I���b6�ӛY�MP-��5�>��J��ejlg�ZF��o&���ݰq!qPS;�AS�$l(�P�GOD�j�c�L�sM��8y��Ư��GA�HwzS�OD�v�\��HK�J�R�"^�~�#c�Zn_����e�W��b�pr�ncq���Ҁ�ǒ�J� �GcO�z9�a�Y3c�M<q��\�N��ږ��gZ����UӁ��Ҩ��K:�0�q�*�z ��q%�{�z5�Hps�mD� =Y��
g*�u�An14��fً�%��#wa�5ȅ��y�'<�_Y��\ߟ��R���Qh��X��7ŜyT@�^+��HY-�L��2���)7���v���n�a���iF��IE2V��t�`��h9��)	�����-�v�.{v��$+@������{"�o���h/��.��k�J���iV��vX��i#�~���F��\�Ĉ�n�0��"��Lt���d��X��K��_���A>��2^{V�(��^�3\�ܠ�r/�l߭�&:���w6%i!fk��9�`��՛��rKF+�W5��m�y��J�ʾ���/lĝ��OJN&x�U��8���>s��zJ��`jo�}z�Vp�w2޺lj�S\굞c����w��^�~��.�Q^��K���f�y:�eV� M=;��D��.����>0_*�U�z_S�_:����u9#xL��Ӹ���*��-(+�0����YI3��6#xj�q"&��&��h��_]&_`�zu���<��?�U��0�L�?�^-�D��KSq�|=�	0+�$���M��"�ל����{u^������v~�x��a��kT���p��`o�_@CNʗ��^ؿ�.�A-�����@g�����0QT�8���Ք��*�ث��E�bm��2K	�r>'N�h`F�����@���D��͗�,���c@-c�Y-3����xޡ7�w":�
�;�2��`�|O� X��nBl n�q�H���e>�Cy�c��su[�Y�����k0#?LJ%fj��	n����ML�J�7b�WljZ^�󥺞�#f�����S8�(}N�V۲ki/K]y����#>>(�^T�a������)qRj����t~z<���;������,\�|6�rۄ��&kE��S71�f�)i��1s�E�^�=:�V7���U����U�_C�4�j�KU+88i����ܦ�\�YIY�z�GeoZw�|CU�[�ԃO�w�t/�`$�jp�FMK0/��,D��v���U�xd��:�3K�jĤ�����>ouk^�^\X.~c:�D��N�E	f�O�����ڱ�d��V��\$Z�uT4n�r�p���m��o�$`ı,�eq ����O��,�m�b!Fݭ�9Z�;����!V'�l�qf�V��1VA�6yD}��p�����Fzsns��ʲ���%d�6��>�= t�Anz��\mn^؁����5�?�7��f�?��u��Yf��q3��JQ䦳)և�9��ʲL�-Y�G�Nk^��x�~6��ڵ����[R��S`��9���#u��|�B�D�~ig��"��Yi�V���B.~%	r���p��F�1����oy��q��j�=�5a�����&���nI\�{��(h�@��˦�C�'�bh0e�u �|�7���[0w��>�8s�a#�}�b��kEB����.e�24��!���ׄ���Qc6�S�Ƈ�'u_;8'!���R�9��E��˧�kv�?���?��N�[�pk@�M��Y���m"^�' �c���-��/�N.ܸ�X�8ʙ���~�OW�Y{� ������$j������Nq���o�>I��=G�%��U�� :�"S�3�G �մ�KQ� =�3�˘E���f�e����u�?��&�#[�&��W�D:����[<��Y��Us���e��"��Lg�=�/��T��_	�6T�7�:e�Gh��N	^�Q,G��!��	�o]��Ӂ�������2C�
��
u��d��$u�X�B�}w��"$ǥ�$�Й���|�W'���SЍ����Y�� ��8�Q�S�R���+�l��Խ5O�O8>cz�8�)l�t����N��$��R8��(vPbNHc��̮���2�&3jnq���R����ӎ+7�osn�J�_� �6mޛj��6X5��eB���zV��mI�c����D���%��8;u6��T*����*�0�r���}W_H~x�����=�\�A���4?zCU��oT�c!�1��#L紺�/x�O���޿��{������Pn�����Bl4�|'��#�e��
qΓ^īIOj�"��L�2�v��m�<�v=n��re	�u�f�81�R��E�ə�Z�zYx�i��>��J.tK���=�T2L8�2�������D3�M�&l�`�{>:�n@��-�"��C+�!�U%B�Y�m�M��aJ��1�eG��XH��elh��p�5s��x�""�@u�w���&�+d��,��cPpo7�c�nBe2��b��6M{�~H�+(���ҘLoL~����Z+�#�$��Fm��W� �X$ �S��HSm�����
�e�!٣Z>2R\,�L��g����˫��W>��^�+��_$�>Q=iD�Ӷ(�'jE0!�L�+]ff�t � �l���4D8����@��^�Q�جޫ>	A��9u�#�JI�k�]��BT(@i#��y�:+�,d�=��<g�y�(f����L��ſ�.�;�9��[&�a�Zǖ:CP"�cuf�f�k�r.&��;�wj-	��y����	'�|kg?���T��@Щ���v�b��p'���8��|�����!��=0�tv�.ϚOx"z��8��C����q�O�E:�Ծ���R�̺Y�OA�� �P{<��b�p���㳹�/Aa��;��F����V���b@u%rc^r|�U�v�)1�nζ��)�-�$����ӻ}f��7|�o?F�.�9i�7*�:�q}�W��t��n� Fb����Gbzo14W��NJ�[����$䀐nQO �Ƴ�h������p(KIk���)�J԰f�Lͣ�%q��>O��R0�_�������6��/q��b��l������4R��V�����KJ/tr�0�OW�!�6�pHKh�V�dб�}S�7�m�ѫ�*��ۧs����^Z��W���<�j�v�,bC%A3W,�sa[�W�X��[��
�OEد��`�������Pޑ�z��;�iX?Su�JZZê3�}�@rX��;���h��vhm��sٗxJ蓮����ڎ7N�����w�c#�/y;L�w]$�8&�?�L�ҬB�9�9���Ɯ�פUO�H ]A.��3n�"���L>��U˥���o�
��G�d*
�]�D��U+&a;�_�a���M�W��_		`�����7n$4����j��O�+�J"J�D%�T��ŵ��dggT�Ѓ��"=H��#��қ�1�iJ[ޝm��Ev��H]�*����6]����Խ8XGV�S���$)���D�jʔ�~�ME�i[��z ��<�!�^������''�p�l<ܶ�&�\h��?A;pp`*L���s��}��c���u׆�`W/�a>��znw��Ң�^9��$t\�y����L����(j�Xcg���Ŭ�g	\~>ÃQ��[�(侾�Pnb��.߹�$�V�>��@�����d��ZטeIX"#�Ą����(��R6H0ZB��$S����yU���p4���z�S�J�����hQ�u�t��k����.���C�|pg���^=��i�Q��%p���Vm�h;&:S�y>��lj������&����o��*���_���j>�ԾYN4��F"Vl���MpXq�a��˛��Q.��y���z�K3���}q!
֪�4�f{u�rݤ8t�WL��JI���Q����w�bҽ���T%_'+�����)�VTU���GHF�5�j#TuDS��Ŵ��#jҊ$��.�.{F�5U��_�>�/����m�
:Kq���A�tH M&c��}蔺K<�|��!	-��K�"=�r� Qq*Rf��f�kM�ߎ$G9��u.��u���v���.R��*|6�
��?d�^%F�Z�D���}Y�[z��kt�>�,L؆�C�g�������U�7L��s|Fs	?�|6����Р9��[��%h�(A7j�]f��-ґx�6�%,lp?x�2r|��)�e�MWh`�����G�ى����_�gU�^�A�i+�B)��$��9���"d��pt�T�b�#��8!�8B�|�ĵ�N���L���jB6��	I�z��h_�`�
Mx�S�=4nCC�'i2ֆ�e�8��D�q�AM�:��+0���h+'sο�b�™mO��	O����Q�ޡ����"z��1�Ӫ�٫Z�_�~��?ϋ�������(Z�+k��eqE��zW���ڣa�@ر�o���U�WO�<Z{�w$T:1/ߥ������ى8��%���M��Hۛe��l��\J�������rs:��j�҈�!.��m�1��[^3�1y�jOӚ�z�������b#��Ȋ��e�zv#r��ضJNR�������9�W���Ϫ��#��!�������$�aD��-�9���S���	�|���؍��F=�!%K�Q�{�x
�zvc���� 
��0��q�r�\�� ?˾p;�~��{��������+�����3צl������*�x S�LA4�c�i:1n����V)�� Z����D ���g�O�c=�Q��ϥ2�}M70�f��>�,��WŚ�	�3X���1ہ�w��'�"���RE
z.��E�J��\��8<&�I;4�1�P¢�-�:hd�F�ݳ��~6�f���h�z퉯m�ܱ�K8�'�mɅE���6���)t���z���_&����3�v���li�N]Vh{������i^�N@v�z�ۋ�M
��8�x}���hB����hY�Nc�U���|�9b��L����`��ٵey`x�~��b̎�uR���뇰�gW,�h�1�^�&�|��K 17e��6���b�|-����&�8ј�"Q�~r�x��mIFEo�:���N���u��Gn7��0�{9Q�k����@7	c.Bo#n�U~�E��@��p���'m�ؑH��|h��@O@,: `�����E/Ӡ�g	O����aپ{��|�`P�+�W8#���:�4�]��A��(����k��*�+9y�gN�v$@jL{��ƺrЄ����_+n����҇I�vW	ʽ7�m����!�d"�$F]q�z	��/��>�u����������_7?XL��y���=�;�9|�H������L?(x�����.D�,��4��4�5P�a2���ݡ�C#@G:��bºFH��[8�3{�A֫C�<��*�D��ƻ��P�e��O̅��~�/:���%���$���Ȯlr�Fy%�*.��M�ы�l����r_��K(���!��/Bz��I2��kFG��l��U��0�k�"޻����~��j�N+�>����1JI����X�n�#���5>e��q+-�E	��N|,te&��O:�<N�&��p8�Z�14{��b偍��G�W�5���� $(�c2��"ߌ��$���������`Be#��֛~6�!.jU�Bě崞*'���/BY�?�&{K�_Ue��^�y�� z4�\�f@�������S���YuY���[�֌:Vqʦc>v1hB?��ⴸ���~�y�X��{Zv��
���L*5V�� gS0���ªy�lD��5W��q�V� ��~��P���ֽf�u���
H��;C��n�x��ȹ������՗$��FM���
S������8�)�υ��sw�K?�׵!e���)�0n���f���қ���U:�pX�9�RԠ[u��MEXO���K�fՑ�h���I7Z�2l��ۙ�L��H�Gؚ�lQ ��x/�����v�8��^��5q����1��߿�+��7j��cE2�8�S�
!�J*d�`Ne�ɡS
���Oͬ��+��YӐ�#��A�x�O����8�8 \k���N۸�Y�,E�qE�<�ᢞ}�_�I��΂��o�r6W�2�Xk(�3/��{�ϧYɎ>�ݾ��t��汀±^�As���E�~��-��ɼp.�(�l�^���4&v�Py�n��ǎ1�9ܮ���t���x$��L���Ҵ>]�gp�?��=������
�#u�U>i���fNbI�Ն"H��m� ��S�cd�!�E�aY���<�n9mv"�N׻"��,�L�D�K���^7����X�Xo�EB],�Ȼ�^�J�Mw�׸�����r� ���k�"z�܃K�:s�1]��pd�j�1v�6z�h�4އAD$��B.|gy��.�I��:�BW}���؟��a|��Uϯ�'�̡$����#���@����\�M����]+\v�3�ᚋ�#!#:�g�cQ�np�U�ۡ���5n�J� �o�r����(�*Gﵢ\G�lF<�s�j�>��v���W벢""�B�P�b�JKK���4{�8�����C��v�.�w!e�B�Z��`���ߓ��gD(�3�g#p��_ĞD=����a*��KyB�����y~�S����r=���K�\4���4�$�mB�p@g�u�6�EfV�]0�Uq���	�7|���q���_�Q��hX��*,��e^'$�W$!~��%}1�?��ncQP�s.���I*�1aWS��n�^�_	���h��郣[���T��|������h���f�nas�mH�8
�=�m���'w����v늊�kr�qg�`+=���$y�OX0��k'\{Z9���V�n��.��w,�`M�Q_Ev��P�ͷs,߼�!H��v�!g�\8�ٝ�)�Jh�\��=�\T�G٦��+xpśe\t&��� ^Z�gw�� ����͛_`��dU<̯C~-� �I�3\>֯��u͒�[�X�$v���ٌ�E+��c�-��~e�4����U��!�E.�I�o���m6�	��A�,_�����:\�ړ���ڰ��<>d�_�R�oU{>p|��%������C��{#�3F�O�p3��/����%'zT���_���ز��'��_G�4������=��wwww��!����;��ŝ�<�w~쏹vg���ꪙ��*��  �7|h����X/K6ٸ���F�7X;��!y�`��v��i{α�c>U �jY+�,B�^ϋk�/�=+���*�6��{�P
��E��{$�P����C�Nے0��v���m���  �0�ٽ�J��a|?o�Gx/f��4S~�h����?0�9�fv��K�kRV�J	N�$8�"��U���CR���L���g����1X�K�C�1`��x��jϽ}�.�q�1��q4w�?^��a�o�x��T\�5gAe%"���F�ʹ�;?�49Uw�	���� ͘�
�$T߉�YY�t9�@u�ĭ�j������׽N�M�� P���<�z6Aj�/�����~W������ˠ�f}�˝$	T΅��Y���?c�q�iMu1�T�<S�*�8e�.tq<&��h�w�v��.%/I� ��۹p'"qk����y�9Q"�1p�u��-J�OV)%��\OR���K�ڕ�����X����o.��k~��:��YU���(�#�{�qԍf�m��A�bMz,c�� {�T����yrܠ_�)�Y�z���2��d�"w�)��Y ��&�����܎%N�74X� ��jƌ@xJ�e�F��N6���U���PU�o��	Pni�qvD9!�͜�[��㰑[8?��@��q��`���g�[��6x>���ڄ~��[D�*-!B�!�jx9�8D$��o۬��u*8�'V�'��-^��l��������sP����m�2r���⟤խ� K���X�p劎� �f����=6�$����0Li���e����'�w��j�C ���=�#�q�&f�&�T��.pO��j�4��U��V��-:G)s�3�oTSta�=:�@����~��=�4ؠo�}�j3i�裛�.L��X ��ק����w���k��O8V�i���/5%c�����q�{KO#
){'�i�/�	�f�E�M$�`W%.��|>��)tz��=�z����Z� @��cgf�����$7?������e�	a�E���a���{׵V�|��CC�qD�>y���7�mfJ̠��8&$Qvg=�G)+�m���x���g<.���P��Z � ����� ��*\�`p�Nh�M���B~����1j�_4�x?T���{����D��b�H�l ��')�,x}�`�9�3���J����mK��6T"*��|�E@s���y/O#�>w*�v	��v�.;'�nT�9�q5��BB��1�{`q��1��A�`������B�-/�A�T�ޓ���T ���wXw8_�_y���|�F���Q���I��+h��ud�5�IAnN�N&T�����n�2 �L���'�iE���B��o��R�����S��)��8�0mRP{9�� ���P)�͇������މ�u���O�L/˃���j9��!�B�)ƸÊ����a�����|�A���6��K!_�q
�:Gc<����� ��	ҹ�����m2��HA���9��/�T9�������b6����������z��q�p·�m��s��C�w�O��/#/� �٢�?S��BhL���Ib�����+h���ݾfg  ��ݐʻ��������6c�3��c��cy�g�����|��I��L�^�C�Cut��@��W�`��Om���~�	po���呋�����_}���oZ�MH:2_q�p@�o�j+�����{�@�ofhm{&ZZQ]]"㺁�.���`$���V��o�Ȁ�.ʵ؉@.��I����=��Iv3:�&�bupO]�\i��^뻼[ߕ��ȱs�;Dph�]�-ǒ���B�;�I���Z�wѤ��֟��h��zZ��&/|/	24���X`��A�#D2��qB��)�g�~�ɰW�����T|���_pm�sE�Q|�X���ɣ�jf�`���ڙ_4�7z-!^{Hf�Y��:�>X����D��:�ύ_��D�A�ۼ��_��Qg�uٽ����~�7��",��U�X���E�}�"Ξ��1�׊bW���'��Thx��;�Ӵ����|�C8R����S�a���Pe&1�څ������2�9<�� ��Ѣy^9l�������a��]3W?>MeG'�PLvv	����3\��k�$�̛���o�ar2"PBj[�A�BPi3�g0�@&�2���3ں��fD&Y� �^���~�yƽrC������ǥ!�I����0h��OF�<�L�6w���g�}_���hG|�D�Ì��_j{΀�����F�n`���B�	l����h�M �0�qjE���x��N!�{ǃ���{/%�����=Z�[�A�zy��`�7��S��'��ö^e��Wyu�.����w�����e'T �2RFo/���Is!���x��d�
�tv���5�9K �y9j<)2�d^I�������g,�P�g�,�����j�5���@p��c��9肉/!#0�A�_����1�\��jq\��i�b-��c�E�b/�!�wdO&S��-~�P�-�����ۂF/e�g�ɒN��Kh#ż<�����j�.h.�;RÀV�-0߷�QZ3�ݚ�����&sn)2o�S\,��'�UO���Îv�Z0
��~ɧ�*���,A��k�[�N���)8O� �\���vc�6����H�[+)W�Fq��ԍDo>�����|��%Z��aR��OakPE#a,4:�jܹ�^$���)LA�t��2�c򈲶�s?0 ta%��i�gF�a�r��I��?�3�����(�W���nb�'�F+���u&�{�a[�<J�b@�u� |��F0OQC����B"�a�=dH�fee�dI���PP|mB��&�}<M�� ��r� �@B�N����@�ps��;nM�D�5���ҟp�?�Y3�R�+���w��b&�4׳�򨫓���[�"��f�?��/���|!"�X��?�s���p�T�\Oռ?��)l�B���,!�5{)}�/D���7���q=�F�<������� n�95Gz|ACmS�ܝ+����a�~���2S��
���J+�r���`�@�'���g3��-%K������T;D�\��l猪i0�Hi��h	S-��Ƀp�~�:�����~sm.��`H�՛Ɠ�(�.B���Էt���6L W[��������d�ĝL5g�a6f���ר�9&���
��/��E��*:%��t���0s85u�19�3[.���?�\�d�ek������j��{U�,��R�əm�Д��3��8�7!�R��j��:�mg���P!ו���(��=Y94,W�}��v�P�?+��GT6!F�!�	O����U�[j.\��|�]/���8�J�5�T&9Q(�ü�+vO���d�H���kE�r.!��wJBRJ���-�͙�н#!��W%�����,�J_�˲��M6*��TX(�@m�o�E}\싕�og"8���&�s�#A�/��SǛ�_�����B��bM����]a��!�{wH����_*�n��w�q-��th0w�ƥ����ZA'��_mf�9�0{�o�_�_r2d�Eme6=�!)��)F��?���7�@c�\�A���y&����f˱UI/n�<��7|��`p0��0°�����_��ί)=��x�X�4�!3�E���s1P���Yv޻~����Wv�C���T~�tJ�)YE��عs�x�k+PVi١�3ڲ�������6ym5wz�~i��>��&�_�|m����|x�laڲ	��?E0�q�rw[����$ht����=6���a�p�w���L�Z�HX�����u�z0N��#1pj`�Y�Gf}�pnEO9�0�����ٻ1��uՏn���+�RC��g�r4 ��_ld��" |�����aaǔ~��I���ۡ�0xꟵؐ���aP6i��%�MMr'i���V��3��ո����5�1��Au��2�T7�+Ͳ�6bkYI�
�#Vj��g�G ղh�w�-I1� 8��<��_�u��ckXp��6�㈉�͞w�W����:r���6a���g:��4$�/o` �H�Շ&L�4������@Oj�T<L@0>J�>���=������e<S��_۱N�:�� $���G/�ְ�$��^-3��&/J��d�z�����  @�fʱ��ߥ��@�k�-��ds5�kG��uU�����"±�&퐥��g���fD��X<(��/���Ĥm��i�W����
JY��a���ґHf���Z��#��݁���t�
~#l�ƒ��#�Ef����=$R���[���8�@���FZDn�4U��̚L���A�g*Ae�����wYDg���r���G��P
b����
�k>�S\0x�0k��V��Y�r0�����
'xUjLM[�5�c-EЛ�wc]�o��Ձ�(9�hF.Y��C
�M<�DLx��\��x:L$YL&iL>�/��Z��C��v���
��Hzh������@ޝ����)#6�7���T9y�~bK^!$���Q\��a��!�49P��nX���_�۰��b��_#�O��L?��ú���I\Hm�r$H��tRk�>�m*������+�r%��ng���S!r$S��8rף��?mq�Q%�{φ���ޫ�|��;{��ȃ�jT��"%}Ӄ(nF6�ڈѐ8瀢J쌸:A�?�Q�_X)�aL����3�"u������
ǳ4YM�}��=�$(�V6��JHj;��D��"c��@RY� ��G%I$=ꌂ��ԥ��m��2��3�v���kCȇ���K�.ɕ>�߬���sKs6R@����x��?T���(v�F����2]హ�������1�l鵖��8�����w��6��,�(HP<����D~���{αÑ���(	@��A]�ܘ�h��Y�dffb��Ęyo]i;��Թ�ӳ�͝��1U����욕�^�RTw��P_�b ���`�;oF񧖘$|||� ������ƿhx��E���Wv�l�7П%̍�z-:����@۸YF���Al���	������f`�'ը�EB7:���?5
��%��*���J3��;���^�{7��9��ѭ`�̄�B�q��T��C�p䝁*/���­�!(�l ��`n�{��c��=�}:4���O���G�ǎ}X�.ڡs�qX�+7lZÄ	b�Ɩ�|�\�[B_u��=����.eh��{�4~{��"����t��xZ�[Cka�SM��g��Y%�Sٴ{��@q0͗�D�$j�}�E5Ȋ�ѠW�?gA��b"����M���7��[��g�\s�+�wdB������U��y9HY�H��r,�Qh�����]�Bbш���qOMǜV�@�opxs3�� �|?��Jy2��9 �P���� ��˘:�����{���zKLF�Ѳ���?��R222�9,�#�۵���kY��ʈp5DHPvE�\��>_5�ө��f�qb�U���T���$V[CEQU�1!ߎr�;\��^!�+��0���`!����	�M�᝭��j)2�Td�A���Ѓq�FE�¢�٥Am~5��ݭR�Z��?�n�Ǹ^WG��߱S@V=D��le+*�x`y����w��.F/9BD��d[����>ǅ�|&vOw/b�s�*�;�:� yG<,"	*�K	Z��ع����n�vT,�h��^(Q~oͬ�ۮOj0!.!j����t�N�Ѭ?�.�f8�1�Po#��E_�R��i1ӭX� �����ٽO}�b4�CBkVQ��&O;���*]g 3��~0�B� ����=�\�:6w����QS����w��@��pxv���C�|GJ\��/�~s5��Q�W�0`z�ðp�3���=k���Ӌ�&��LlG@��/�XLydoE�FR�-S#����q��-��̼?{7t�U���i�z�u��@��
�af���OF��{~^�	bN_qw�z�,���D;��܇q�x�4�G�D�����Gx�2V2��> %v_. It�~�҈ڪCK ���R��y~N~?�s��H���?�n��_a�dK�����G^�� ;>mc.�����h�SiuWe(�������\x�����1(��,|��(!���}��0�:q䪆L�9�̆^L_�����_r�����A�j,*t����m-�!U�R����F0p���*k hZ��Ҥc+p��BH��u�~8nr��oop�غ�<��|Y��jqq/��׬a�J��<��$�_�Sh(]���]p��Ad{��(u(?#���8��K�Mx�I��y}��M��q}0���5���H�{�Y춗a���:[=f��	���ͳ!s���Gܢ�b�!�as�2�"cP`h��rL���gc�Y�p*���v�r�˷�_SZ��2����L�_̑�gJ�*���S�סU(o���� G@-�5H=���jNvo����ʼ֣H�]T�]�&��O2�/��Őh�(6w5O�Qm�����&�(\��Nx��/>�9^�p�y�H*L�9ge7���8���杹WKoE���<6G�4�	�ٳd�u�:�8��ݐW��9ˁ���M�S�j�'���7w��P���;�so�S��JgI�.��3<��gً��;�~�I5��X�.�����*!�s��,�)�D����7��w�z����_�)�ɤ��wR�3s,{j	�4��Q�ĸ����#���|��~�G�+V�����3F���� m�'���
pi/��VX4�+0�@-� ��뭪������N���˜JQU�j+�a�X=����<����.H�aI��ʩ���i��TL��4b�}� �TߝW_Q6��L�t�Q�\Ž%���N�aҏh7t���@`�D��k �Rth�`h��4�L�m�G�#�w��_�{t;�Õ�m�ʚ�� ��ؽmu!��|�$���h�V�i�a�]n�j$9W
�Ƣ;�3��xWloG3ZI� }c�,e�6c��0W�,�����P�����Hdǧ��m\������M�I�m&���C3�͎�F��������f�M
�E�y��bL��K��`Iơ����a�$FZZ�6`� C��f�j`ъ��s��~�ֆX��ψD]��/z��H�8���W�Px�Q�t�u��e7%�m8?$�vY��1g1b��b���9+�/��m�4�D
P��藜����A������F\`vx�j�w`�&�Ӣ��lQ'}��t6T?9� �o����+��$��Ck��"�\�퐚���得aV�y'Cd�=�s���*䥭&�.NOEyɑIW#�6�/6�De�B%nf	�oX��:�&g:��> �[�k��S��`���܁���G�`���!*�c�+ȕ`ߵ:�ff}�6��ұS�iuv�m|�16և�Q^�6=^�"W5v��Ԉ����5��o8<l���,��Z����ֳݶ��Z���,�e�VSs���Gf��@�zf.�d4+Ks�\9���CڴMPh��IWۖ�tZ+�+L<g�s&�^��_��
!�=��n���y#����J�d{#7�ע�R'�z=���E4m3m���y���׌����3RhG���i=-��&(�����t�3����AuJ�u�4�q�8���8��A�Œ�L�n	�*\'�������%���Z��r�wm�� m�Ø���{�ع!�c�H�~�ϲolx�9����ld������5�jb� ��X1�H�Y���54hH�Sۙ �r����ã��Q�2��KH��7K�=��5��S��V��w$�����8��	���?���=3�1��{;�U�#!JJ�a�G���ȉ��#>�h)Y��oD��y0F+��o���֕���0�-��o�O&�`��l�����l�ę�mHI(p�U2������� ���ps�RĸU��!�י�i����aZ@���C@��\����ɕ�
�5�a�B
4d�Hlr�������95����n���V�I�P%��[=���f):�lS�/,p0���r�{<��?OL����!Rݞ����V�_/�ea������ެL��v�v��~��E������P�s��&�����:�����%W� �-�(���<�l3Q��Qf�~�-u�^����٬5p��H�1��;�EZ5'�r_�'2�.d( l��A���H���y�iø�$�M�_gq>F>��bܟX�9��:f���E�,oy���P�����FYL��Z�fo��Eki�]�]�����F͍�Q��x�w�<}Դ����o}nGAt`P�S���E=���Ǹo��8��}��Af5��mw���Ia�jW�{f��fkL�
�b�
"�Ki�u��s\���S�n���x@��uw�� b3��)tM��x���VS��󭏟��d�,ǵ����RI��J[�i1�/��o�\�R�7l��
g�o2�8q����la��m��r�s!�2�:���,@��x�M�ZH㯀Ͱj?+n��̎e��u�x
�!�fE�^����V@���.�K��
!��ԋҼc[�)<Ͼ�`�����n���of�=��e#�8`�O�%��'��������7��b_��D"~�0J�gp��R�����\[,˘�T�������m�7'�_�i�UB	�U�^Aj�;�!E/:h��S����{v�m�v���lz0��i~��=�YO��x��4�އ���3�ǽ%�&�c���
�g9Ӊ0cŗ6����}�A�$�#n��I-�p[�� d�)���u!��b���?[��r�T�����:�	h�^h�b�I����_g��<��e46B���u�>��cv�L��a�]��Zm8�3q�N��.����1$���6��5�%�K�jV�\f96��b<�?с�T�_�in�r���3�s�q��1�1$S%_T�������J1-n&љ�d&q2rU�o���Y�W�.���qqɥ3������V"�<�=���NM΃��Ԝ͑N��e�4�������X@�	�����6N'˧Cf��fj�6X�dѮ4��͸��f��j�I>XB��y_�O�}�^�!U����DC珌�	,ܤ�y�It���su���(��j�� j�b4D��Y�f��*�Ֆ�_x(sF�:h4�4x9���
:<��lZ������0��[H`+���l^ѹ<��F�8����o������:D��vZ��yI�it�;[0a��A^B��|��_��7�&��/F�T��A78"C�_0ղ���N�{*��n�e�
,ڰ����-�t�����j� ��o��_J��n��E�"��lM,�]ߖirl�3!c��*~�9=I�e`	K��C�R*3ۊ��pm*a�1ی�{(������*Wc�_��[���)�c8������0c}��6Bf8�~�JJz��������Tb75���!�_q��$V)���?���y��D�ww:��{-e8�iru�K�F/�aŎl�|z%%rm��Î)g����4��@���P�XjO��^89�I�5;�t�����s�������xŜצ���uC�g6\�hh�.�V_1[U��q�����=���9�|�0WX�[bL��mC?�47�z��ּ�|���.���ְi0`^���dG�����P֖k�;n��.��|�vm.�ĺ8�MM�/�]�q��yO�^Y�1U���̳�`r�ጓ19�RN>�Y��)0X(t6�.��S�X|�l1��a�[��P8�q��q ��u��^�������p�"u�/B�I��:�v���1��}�7��7�	5qg*X�80^��n�,��pP`���q����l���l:�,w��BPϱz%5��_���������~-���Mc�)kf&B�Ÿo>Ų��LF�5ε����Um�"�B�g\��7QA4ؾ��q�����1�56�ɴm�Co�7禲>�E�s��v]I�
;�VE]����x��p(�sV ����ju�C_��N���@/N�}��`D��:C�".C/k�����}?�wz��ﻥ�l�����h}���tR;h����"��]��UU�C>S���kx�_�O�X�	�K�T$�tmf>�ח�տ��g��+�$%d��jO��b���#~*�WӋȺ)�B �9�+�c0�B����7O<I���IGX��x`��0B����s�[�"L~�IN(:�v[��n��,Q��A�ׄ�z?��� H�S����WWz\U��n3������<�:-�@gY�M�pC�J,��rs�'�O���y�?;�3�Lu3��i��(��U��F��g���c�0�x%x�W���c�dC��b+6��M��Tg)�)���E1�X֦��",�e"{9��6�K����A�H�u�P}��x�1�[�<~�GBϮZ��k,�oŠtk"�Yǒ�ޖ?���r]]=�&�_*�A#����Q)�;v�6�@����Z�;��\��}E��C��{u@�^��J�2��SL����19�i,:�	��P�*��<pU�1r��Z�n�F-�Qv��z�B^��δ7;�(Ӄ�(�TF��?FȨeV�[_�7)�wY��Uݗ��Ӝb]��w�����y���C������$�?k�o5[���^3�:������®���t������l�g�f��bu���%�2r:.�Ű
������I���_��^<�ü�=�Eo�wK�hh`�måC�W�~،&u6=Ԅ�^(�|�~?jo��ٯ�Y�W�	ِ��Gy��?���霁W�h�!��(Ѻ�2n7IR(V�@2�?e�s�Af� ��Vy]�=͎�I۴�J�7x�X���L6���F�!m��b��bm�X_��P���D�bN
�B]�kQjyNi�_*M�Q�r���\�dA"��Q-"*`��e{p�s�rcv�=u���>��O��)Ct(Tz�����BKA����\���$��R�6�>��Kq�xHmU
oy$��kd����0��q�ՊdQ���ߢ)H�2�!`�B:A��Q2���K	�{��},�-D�^Xo�#���l��k��{��xkl=�6������<T���t�N��cgt��o��� iI��qs�
���Lгk�e��-�T� ���lԺ��dڌ��}(����1�f��fq�6szq�����o��Ǫ�� ��O�ya���ݢy(�X𖕆j��+f�;��?���]P�17�d[q0$�ѡ  �HB�?T�Bcks�p$��^�BYX���P/��}�@�\�1����]$Ȗ&!��>��P�݂��4��΃-t_^�G��e�w���bŜ؊�q}"bVl�M^]?^��a'��a~Z��)G�z����E?��Xq�.`E��VD#!��oo~��c:(W�n�D�C�n(���l$�t؏��l�H �vB�2E���}��~����y��p��Vk���&����ުb5Ͼ����+��D�]����0��G��ķ&�r��q�`�js�n�p���%��M�C)=H�0k�o��+�Q�H������Wjм�4bY��4~װg�N[�����0U�R}��RE�I��-�kP��C�'h�U���>��ו}��I/i��o����7��?k���U�?5�'و4�Y�
b�\<t��~!��WPss��]�!:�2VjV:�O������(�A�uM���]{,��^��H]8��g͙۴�0�A#�at���e hĝ|)�Aa1����/���xŠ�V-��\�g#�e��� ~���_x����AU�1��ɍ�I	���b)�[�|W������.�Z<�8��9�2�{�?w'�ɿ��:(��s���!����A�?�k�����}��J����:�x
ʛ��S5X$fg��uB���!�����t*K�n��l�d�sq�K�]�/8ͽ��Ƃ�����O_�(��K;�s��s�/�%f?�YK?�,��D5�:�tnlO��G�6{y���s�В�rt=���u�= $CËHi,��"d�zit7���FR����ۜ����ƿ+';�H�T.���tj�H]q� }�����
�I��1�}#���<]TK��P4K<w�Fh�9�<�&h�x��].����'ep���ft�GQ� ������q�^�k/���$k	�!�$�
�M*���ɨ>�wē�G�-�p���`�4T�̡ydwf�����kU���W������s�i��|RTf��LR �<t�&�	/��mpB]f�9v��(�7�r�J�H9�SIom�ˎsEp��$�䒊1g&�f������F��c�]�ujP�LXq�Y{LA֘/��d� �K�����NgV=3ʺ�u�N~C���/������2΋�K��[�:k1�8t�n#��+d@���0z?�>H�����YU;ѽ�f�Q/JH���{=V,�����v�6H���b^������d�|I
��ԛ��tgj�|�Gl��m�"�o��&�_]������BGz�s��cr�	IEZ���fJ�E�1"W���	)KZL�!�Jm���;0勨����gGu�L}X��I��Qf��I2��ӯ�lI��,qU�n2 	�[���8�7~z�1�3����wZo�G��$�1W2����~9�6F�������M�9�Lyht|�T�lpr�R���2C+��I��r�w���_m_ig�Z$�%�2��TX�ʉR4�;F�wq�~�>�5��-��D7����U�P��٘�I�D_��Vi�]�;A�����n�5��т-"����v`
�\j+Q9W����h�D�
����{.L_uBuN�#���xhma��>t��ҍ`�v�jI]Ex�p}DL�í?����Z��n�&$B��CD3�%҉����A�Y��Ms����5�0&B� �~�O�wP��8��Gg@��kY��0ƈ�+H�7�Ք4Rf�He��!��	����>C@��c+kѲ�(;�$��Hp�h�4��D�_�nN��E��hX�S���~ڻ�������y4�˾:���zY�8��.���gt3��,E^!��e����`hŊ���ى�E�W���,��E�e���X�$�> ���$�&��]��]t�ߎJ#@�� ��� 0Psގz-���_px�L��V�K�u@L�l����k��)�Ԡ�-���+�{�c�Ѷ����,���x�di8�p�Z.��aθ#	1Xɬ��	+��mX����󯾬̾}��1:�s�~V�x�4K<I8Wg�s���R32Fܔ>��U0��Փ�)�-��o��������M�/�̵�TJ(ע���9��H$=�j�W�,%yK�3��ã�FƆ����p�������D��a�uy�UB�r�_�d�����N��
��tE�i����$�#ǲ��hq�C��L|ű��x#�¸H<�b�/��;�i�@6M^��]�e_�)�x�I_ڮ/���}�`/�����R1���Xs����W��8_EO�x$N2��P�:(d�ϻ�W|ْ�xA3
]Q�j��<��[*�ȧ�PjNA4���.T�=q�]w�%��<��o��A]I�J��m�p��7��n�pO��L����IWoF�}�y`�l�Ӏ6����̄�q�D���`>�/A}Q��$A|"k�����y�]�~�I3�|O]#���yI�y2�EI1���/�7����Y��	����@'q�zY��K7)�����d�T(��7Sn�������E��ӓ}B��8�J�$:�O*���/5��L���8;S�nn�0�}��.6B�$��7���/)�� ���ȠW��o2������u-}/�t�����c��f��8G��x��$Ӽ�恮�����N��6i��D��y7Gui2�c�>g~q�rwJ���T�@��v0�lE)�ビ>Y�����h:,YF��Y6ܣ��0"y�*Չ&�m�sX���P�p����n�i%q�����LE�XW�23�w��^s���e!Lb|i�]�'�X%���� ��G��'Py�4��7��	����`��@�����]F�)��p���<�wI2�n�����j��wB�I����6<��V�1�D4�v��D��&�7Β�f�(����'(t�/�,��WM���G�U������A���p���w��<|��jbH��2�:{J�"I+nI���p�m���B�����z��r�PpQL����Kj��̨��̢��M�6��G����"Dp�������%��rI~o�T�1�(x��$l(Ƞ���=�c{5 ��h~��)8��.ie������e�%���=,m��z�l5����E�؈t2 ��'�A� ��$� �=��L(��^�Ϲc�J��)9t���8��\��oV��-��B��%p.MW��@��Jc��ŦZm�u��Mu�,j�0N�UO�JޯY��{��3�3��)1�����!5끕2{��e�P�MA�5���� 'Q��z���##~e�+�O+���w� ���X��f���PZ6L���i{Z7~�ï���Su��-l` ���5�{t�k��%�ز]�zVJA ��~�Nt���V�!tVa��Mj���jڬ��)-ad���Z�)&ą��͔�8C�*_�x�z��m�����&�?�4I�W�|7�!T�.��g;ڗ���t��(A³�_E3�aqΈr������@���{�Y(M��b%"�\|A?�	��y�cM��(C�����%*�ϚhE������o�Bvm@��~,�q$l�?4$�|��V�|Ջ�sB[��0�*.�
�>X`�|p��l9M��X���c�z ��Ei��:���?�!��ST`՛����z�H�T#wK��|cYE���;�n�ss�jLtk�8Ocz���G�F*�C�m��N\B�)�n����R��y�n�%��[W�y~�~�I�(�����Z��k%:%]�ڷA^C,���E����vO����آ߈'3m��� �@?�h~._h|�����`�c5H�0V�BÙ������0�Ϻ�9�tNf3�^Ur�L���ϟu#�)&��ŀ��VgZ�O�#�F�('�E��g��
sD�G� ��i��`';�~�J���ήb(H�V#�Tw�y�x`/�K�86	��m�'����qZ��֭�0������3�C��cSi=z�W���:����6��|9�,�Z|�r!�=�tX��Q�0������y!=�85��a�c�ܺ�YSAz�x�搫e`���Wj�p
��+3��j��	��㣞[���g�R����Jn�,b�a6.(Ļ���ފ��ԯ�l4puT<��KF�U�s��ɫ��� ����,yۤ�^��1"�"����V�*k�߽��E|a-�@�Ƶ/L�zW�,�tQΥ�KޱeYa�w��i��gr:�Z������N͵ҟ�j�:>c����h����:G�����?��4�=G5f���<|�&} _��Q����ڥvR��8����u�ƚ�ԲK�
��0�� f����:q9@���z����߫�^��~kI5-�
I�J��X�Nj�w�t�>�w����F�6�82~�V�ۉ-;H������!�K.��H�f��<6sh$%��๜��q`r�+f[���>��a~z���]U?�<�ql��EЖS2_�h�thR{Hv�,*������*���|tj�Ŷ��nemZXɣ�?���ƌ��p��B��0��,�3��BG�����Jx1��b�=�I+h����Ƭw�Nc��>]m�|n�����f�Sg|!�Nb�h�mC���I��EX�gz|l������p礫e�z������{N��]�����e��׌�|Q�.�����&�ނF&��26�� ���q�٢r���1�w�yS�R�(-�8�����x���ز�ym?< Uxҋ��_��䂴wb�ԫ"Uy鋸�eI���f�U�O���wt��se7��v�M��vFd�2D���z��gV�Z��s]��=�E���s����D\�{v6u���-�Uἑ���z���=�9�����ɂ8:\�>���݊�j�ө
����0��Ӗ`��/7Z�v�F�es�{�\p�1�� �q��R�����`5���v�mڒ^���c�L:���C�6�)��!�3k�aSr���ý�e�O�	RX�/�f�Նۍ0����k�+�D���(_�ˋ�c�0���-0uE�V�m败����#8Xk-�w��J�[^#�U�NX�I��-��u�?��4S���fN(�:<��݈^���5k��T�Ң�zf��R���� ˬHp�`�"X@�N�x|L*!��ȳ���o�r��4h��&+�BgJ,��@S��	մ�܋Z�����W;����ռ;W슛�Vj7�Ȟ��2��-�&���ͧh	+�� �2�MlNw��̿-��.��ë��鉶t;��Z�9���=\��fN�ܚsJ�%����Y�u�=\iy�n�,TFW��z��W�JM�T�Q�i2����g����Mt��jl뼬� �?��(�`���@n��!@��%����!�;�����%�����7����������:�w�^{�>�NCR��1�[�����}mF�X"�#��/�d(�[�S�!;s�{|��\�#��N�0F}7봥C�\������R���`x�n9F�=1��?��J�B�r+Yº����Dֺ��_�i�.�>��SV^}`�Ti���W#=S��FV-�Q��D$��==k�%�bֻ�\�?����р�_f��'e���*����{>b��W��t��K/�ڠ��p���K�էm��"�B+��4����&%�����M�_�l^K�Xi܎>�]o>���D���1E2n�9h���~��)"�4�������G{��.&Ib�-{{R!���bR�Uv}�e�q�Gg�$�Wj^쑞&��܍s��e�LP�Thl��^���u��<��o�k���^�/� ��ڐA��/�3c`#����rh:���j>���X��k�]f!�xL��o���\�	
�N/��ܓ�:������;'|Y��IS�[�d�v�3M�9�G�oeD�0!=`UT��c�˺$0���[�Q�b�\k~�ᏸ P�'���HeO�3��i�Su��8�lm�k����)��e*l<�,Ⱥ_,g��:T�fx�C;ק'���
�6��U�]��n}h�B�<'���pS���g�_�.g=�����D	�%um������I�y��uE�}uZ���g���&�-��n #su� ���/�>8��Q�q�-�_�_���f���=t�[�2�[���� ��&F݉L�	�s�˥#�g������zY��o���ˠVf�B���Xq0{hge� ��m׌���s\;#�e��ʺ���E��=�����fʟ-R���e�	m�3)��q�=���fT�~�~+�o:���?B҈5����^��tKy�چ�}��	KM���� 8�i)Ŏ{n%�����s�
ZQ�>b\�B�Y��I[r^�M��v̽����z������q�\�&>�*�{���|�bA���w�nX��#D��x�����#��	!���JB�O6'u�?�v�ig��m z��M�tD;{��_���B���c�����^��8RF�6�"��������$�k/������V���۾��}�� �D5�	CU�;�o�x4j_��e�2	X����5�5]Q]%����l$.m��7?z�Jj����}׬�5��
��a����v���G�]�y1޸oK�O�!�d���iY []N
����QlYa}R�_��Z�L��2�k�x���w�#9�'� k\�w3�R�����hK}�۟�)~	���,�|�FT���&�z�Ry�����՜��r��
?>n��^Vtٲdm��>� ~-�N�C����$=À��M��f�S<d�Omac��j��H���!me�E����(3�����iǷ[.�	�iD,�WX��'�7P���k�MK3�i]�Z�|��m�qU��$I�x5)�G(9(�v�W���Ⱦ���S�
	}�Xȱ�ѪO_���(�e����SBi�Q��K��*~�pd��)*r4@
��%��_�� Q��@p����ӕE��|;�����6*3�^I%K�]���J��@@��?Κ���a?k�1��gǃj����Z�����/�)���v��Θ@*X����)�a8�4���Qȕ�����c�r�}�sm)�e����h��NT wv�Q�:��!�O���P��BߣT������K��A�< �e�����mmE�s�| m)��+�������K�B}��Ɍ*��3�.�k�8��k�U��i~DС��['�|�Ԭ��ur����f�����=
�W+���k!�W�����2߼���?\c�����J����~��j���m�}u�����y����lfJ�p��:$��W���������+Ǣ�L&�k������:�����0=�̦��X��E�"��B���s>�<crFӹ���7b����r��/.��3M�l�~�}����+qD�Jڋ^[d���W�cώOK+�.�0���=��mj	x���4,��*����P�8������L�{^&ۇ�b<�E;�9��XsF�e�����˙hĥ���CWB�8T� +9��O���G=����չv$�N`��*��"X�bC���Ҏ`�ި�b|bʵo�50���D���T�GrZk�qa>g�����mx5�gJ�eI����T`L��]L�D �$q�9���V]�1�.H��Ի,a��T���j�?ڭ�_<��h�9-#����0��nE38Zv�PZ��P�GU�f\��vx�@f��S��\ѓ]�ˈ�ÎW#{R7ɘX[.��T�!���ʺ�1����q_�IkRg��M�_�f��K����$��,\��ևhh�o@�u��S��rq
���}�0L^t�	���H�緒��9T`��x��aߦ�T��p��fR��/�bEf��a)w�V������ntf>�IF��ʑ\ӄ�vϯ���TVjT����d�S������
��e�i��y�@�EA{��w��T�YG�3�h�p�E�i�n�ӌ�o��eB��G�@S���w7�3��,|�=���o�4��e/x�%��
Z�٫�Um$?F�����L��]^s:C�Ϥ�3�n��T�őh���~�r?~*Ֆ�W�h��<Ϯ1�c�`j��Y�����-�[�o�G��OUZ������kL'���h�u��H�r�u<>�c��)fijTk��.гP�Y�u�14��Fz�F�٥�ͨ�[+��7PY	p���d!%T[�����/Np"���Q_s����|�~)��L`�/]_8@9ؕj_����K7�w��N�(Em�Oc��^�T�8����� X�=hVBΆ[eY[)��\�)��$���܀(_{B�;�w5�G�{�Q5'eb:%L;�hG+�l ��U�35�6��؆�KX����EC�m������( C��9k^=���u���;�3� w��T��Z�ph9�cu�#�ԡ�f���f����������l���lɽ�<����L1I�ǉN$�\e��,�jӵ:2���~��۳:W�E�m��2�OCӉ'LH��!	�*�a�/d��i��̫6�g���<�1~����YQ\wU�s�GQ��2���U���oKA1����ˢ��u�}��=$��K
o�lZn[ �\z��XA5F���g#V�	���E�e��쯝}(Y5\��)X�A��+�P'Q�)>�%�o�S����?�͍6fĩ��x�m��y�l����8��f_A�w4I|p�XL�	��~�p�񷧪��3�8g��'5���qܴk�p�}
�^X}N7�+����ͅ��=�I�T�jl��f� ���֡fL�M.��Ҡ^���1�L
x޳���s��/kF�����4�3DXe�8�V�l�0JyfL�J�|̻�8�F��^C���84#)����X�?�\��H���؈A��&�3c�Dfȝ�w�[��؝F.��it#���2ԧ3q�z��6��'/�7>�zʱ�����$�zH��P4<���	a@��K�KMp_wl3c=L�Ģ��Ab�y*]��0�B0G� έ�z\:Ӫ[�\S�	�C�DH94r6����P;c��z�O��F�����uf��âp.*VM�u!�ѽ�Z~�j`G���{w�_����!�Q�iX�LդU\c/<�+�XA#�a���D�FO%��.B`֢!Sc"�)���' ���׽������s�:Fd��s%|]>|]��eZ�zq���5�_�Mh�kpi�I�rV͖U�i؉��μ
���b�-ϱ��[���=QEB���u1����oH� :���9�
a�&F�/�/��e��;�`w�����w��6 �*c%Nh7���y=Ȭ�Ǳ��Y�Z���f��n�呒�޿G]���`	#f��BL�����ȫO��ߪ��?�%��Um0z��Q�Z`�ƾL�p�7���Fr��M��Ѿ���T�& ��G���;(�u��xq�~H��_�+��[����#���gtÙ��;
2p'�E�%��1��� &�X�g�&RK*�����t~�"�7d�����W��>�m݌}�nM���%s� ��Lim\��A�p�>~���+����d+}{텣a�:[rM#v}�	�1�!�Ew�(Y�Y�4D�Ƕ2�DJ��9r�<F�W��P`�wMs��{���>�G��/�Q��|:�+M��fQ���'歝}�W����Q.�s,bo�Q�g#���O��:���4�f:��v��bfL(�������˥�V�Hwg�x������K[�u5�+��o��1^�>�0���"c '%7/���Mi�"Uo���
�\��� ���Q�/����������TΚG#���(���?f0��qc.�/ �!�����H�C��VU|��E;��FE��4�tD�A�7��E%΃��
�g�*���iqs�3!.;γ�	"/pW��=]�=r4��!����.�k��D
�~�e5����8g�;?�x�U��~ҫn�N{5Ƈ�1��@(�yX�F�ү�����~4~�T+��+!9���N����
>��`������-1�WƘ#UJ��������"sGES�7n����ڡuX҂{D�S,?+�a����^�X#	�; 8���;lDF��ɋ�����`�ͤ�*�2VP0=�����
��^�d�>ݒ�l�W{m��@�v&0z��!L�*�I��w
�P�ϔ��Ә��U�	�O�;T?�/l����[Y6�}�k�]��%"���Ũ���ހ]�N�]�n|B�vk#�b�cMy�A;��*�s���e��/��:� ���q*ސ������/���<T�[��J�i������2$��V�Jۨ'.ы5 8|�8����u��5�!acb2 |$C1�plW��خ?j�|O"�=.?0�����0j��u�fFr͎�|�p�Ci����j-�Y��u�d7�Pcp�c�G�9:����A屈r���*�&@EҋK�DWgrq�:���H�3��q�a;�����u񲀛��&<sS��=����4mI���ڻ����ߞ=������s���z�dm!��6x��_Ҥųr���?mD��Lh�C��MZa��dZ�3���:�)#9V���~��r)�_\Ǎ�]�]8Tt#7�Q�y��g�0K�f����g�XK>|�[�9_s�7����yO��T�?�+�)@�[j4,�;���r��L�M|?�B-:�b���?�~�z++	A���|u�R����rԂ����V\���Gx��H\�}���|� 6N����pV�z�:�<�
�V��Ņ����!X2"�9t.������m߇d�:���?��*d!�B��'0i�Y���w�TaD�3M�lk����,��Q~Ϳy��t=J����,�� u���-��j8�
�1�f�
��żf�0}d���U,\Ij����H��3��_�]���Lѧ3�"����Ɠ�nuz
-�C�/��������}Aȱ&ɥ��;:T�wq�%��<6�2d����3�n#�Z��y��̝8���1<R�)*a��s��:1�EU�����ϖ'b�:���P*�e@G��a�3�@������_N�RSU,�~U�}��8�Af҆�tJI�動
R�dZ!v��6�o��#�v�������2b�<M����9�����jئ�d�R����y��,�����@�D+��~w�)���a[t�I��::���g�r�6�_Xd,�?x=�q��f��~�I^#p#,��6O���-���=�^|���g}����,�-�^�r��#�T����.����E���5٢�8H��E�Nl
w���VC,.������ *�����A���`��R�xy#ϪT�mW�`�,h̤����GOko�8����<�7�����b�0ɋ�6�'�]|NIT
�wgұ1A�x������fnu
��4��BX$�,��Y�Q]U#�����c������_����㸗����X����n�(����Ǣ6M2m�A0������<iHN`�D^H"b5�5��~"Q�ܨ���E���@�J�T�S_��O�/w/kA�.C�c8�0�P~��x��$ICma�� hV�2�^]Piĸ�we� 4�o�os��S�S��9e�e�=^�"���qõ�UM�{�1[V����%$=�x	��A	Ұw�]I�S���!<0�*����A�O����A�`��4�O�=�Yݏ��sڪ�ά����_�ua(��:�"�����C�~s|���V*4�W����H����JRK����&����B�5C� �կ_W� �8z�፦�2f$��kj�wV1���p�v����k��5hn;�b����sڮ�u2�%?��SQ��JUL��0�vHd�P��ٺ�����4S	vJ�.Q�rX�L3-EtG�t� ���X�ӓc11T�b�*��/p���H�O����7���L&�L'����2�1�f��Hd)�$�<�z3#k�ȩ�$3�}P2mX���0�f����⽴ng�NȠZH���;5M�L�lmɅ��C���U�:�M���ȤgEzp��݈�����[���Y�4!��U�T(�Ĵ$mt	EQȭմn����/����B�H"Dޟ�ì%/r����Y����_7O�Fl�~N%ؖp���Ƿ����$]�<�7�6����˙�m�^���"X�O �c{�������gd�~R~��6�{�16ق(�K\��9�8!�������+��)k�ˤ"
�8US D.���w��Wo.�x��	P�/��J�B=��I�0�Z\��{��A��O���c.�Y��I�Xj�kT0�k��< C�&EVU��fZ�:¸��G���P� w��7>�D��|L�m~��̱�<��P�v��6m|O�G��(�Tl�^!R_��W���_���\�䣜���3jDHB�$�W�)X"\'3 Q��o�g�� au�T�)X�n��T�:�`)@`�+cs+T��X��,�0bf8\f*\p��Y��4+!�� ӳ��kt���H�Š$��W������&TB�Z§[��������`�cdGB'!9�2�2��[����h�?>C�e�O�~�4�F{v�8O�Ma�}2�L��l�G�'��	��{�����7��?F�%�!:�.#L�i�.6�1v�������X�P��!n��"]�	��?��,�D��=\"����E��čMDs�D���b8��b���8�,���DK6n�����9ww�-�x��uT**>`,fW%b��5Ɋ@�
O��W�[�j���^;>�Ҝ�)�_l�%{A��O\Z1�FD*!�##�|�|Is1�rxsm�_�����Jۓ:�ۢu��N�A4�h�)��B���(�Q؜�^��Ԥ��r�RA�|�zJJ~5�-���ϓU��'�v�,Ï}<�[��i���'.��Q
��
��3���\Is��k�k����_��U\x9~���I�w���M�q�v�	�A�Z�3��G�k�!Z�����*�7J�	JqX�%����(�Q�z�7�����۴��G�	!�C;72���Z��#w���z�D���S��ng��,540��:���!�������}�.�k�S�?���q:=����������E���UnRv�A�Q�����կ:~c���<�嬢��{��@l�|���h�~V�Z �w�s�
T�/O�l�4&b�0M5)��x�d�ܸ�6#�t����k$*.�c��C2���TN���Eo?bq��ECuzc��3"�hţC���(�+Wz��@)�06�8e �|�CR.�v�H���9��KPT�8�߹�����3"�.Lm�uuxr�ؐr04$���԰�('+Y���?��'(�Hpk��n�����!�ed��<V��JT����NLl0�5-�Ễ扝���"�_VE�	u{]���?�>5m��j�ҾOP��s�ʢ%*y��@-�5�`��z�|® �Z��'�r�;��OVH�_:�����Bz]�XyڣK��~�EI[��tJ������H�o/���ƒ���k������|�������e��~�J"��hj�*E�q����)�U��2������ƌ�i��%Z*pvV-y�c�M;��yW�@tq�����n��?�:�������<�����t..;������;Ƚ/�@�������Y��E����PK�����?v�]Qb/���U[<�{������$`\MJA���J��vv3�G#H��� à�Cdbbb&ՇDHwm  a��?����-j��4�f,�#�?f/&3���6���ۉ�pI��PD� %˄�n���'��3O�'�vcк�r�%`/(��s-�)�:�K�F�T���`�#�5(	I B����:�[�
ނ����be[{MC�m]3����_�F:�� L��(����E)�W^�X�[�-�B�1ۯ���? �3zUס�?�_e���+E�#�MX�#�F�6M��<+¥t�0�v~xյ�`(�J%Įa�苎1�!�/��D�"I$����]vJ����\���`��m���{Y�g��m\��0���R�(�
�"�֐=)�_�~}i��ߍB�T�%�fMKT;�����3�lz���Т'�b!IW�Ioe�� n=vӿ�;�kS�f�c�n�K=�^�+�Bi�~ѓBTE8�����4Т\"!&��}k
�7�Qu|��?Ҧ�	���v�c�t�	L
0��N��F�����
�E��L/��Z��[�]�e��k���	����.�����KX=��+�6,.�ЩMp�:i�A�A )�K������}v]�mD2sq\:�J rt�8����l��@�O�Դo����6GV1�F�}n*�դ(��D��4/��]=�%qcʻ-���f�Fb��ۧ��c�	o։�}����=V���&�_p<�OA:��U���yF�v'������K��y��W��0�Ub�R�XMhﷲ�������|�����J2�%yF(�_cDj3�n�m��1<���<?�O�8ΟpO*e7ѸR�C��;�	x*uE���,��>���ǯO��CLΉ��t�p�?���0���������tt�'ͧgf�F�~��(2��-�n��0Ǯ���*�QJ]����8��@��."@��-o.+�蟼uO��kz,(�j��jC�:�c�#���G���� �m��<5���B���b_�f���Up���c"9l�e���O9բ��#�oy�TԊ;W�X�a����.��2���o7�Ј��׸���N��[*)5\� "&���;�i��䱆����?*@�R@�騈���.X�A{���"Ыߏ���%��P8^,E�ӫ�P�1�<I��7��.:���@�IVW�����:K)�ķ&$���#j��A_�G�ǔ������5c����0�ｑ�j��t	8����\K��.u���:���y���>b\1����Jߊ%�Z��ƾ�<_l`^h�<t���~�"aV_�B�/l[��vj"��[�^uʺ�����iD�������eRE�:1QK�'�:���ܸR�-,,D��~���C�5Kܺ<�g�̸�{����ʠm�̇us�E�q�c&�\�/E�A��`�m��.����_�P2�?��Mo��s��X��F�X�9M�RQ�%�X��Bz<E"HIe%b"�ԲRy�����*�㨄�<Z�3���Ȇ<�~O	�'�@��	�^KjZ��ii�Rﭝ���띢H��N��'R�e� /�!`��$KÊt�m����l_V��S�Y�6t����@�a�Z,kj_R]xm������eo\��w����<.��Yt�AN��W�9�Jk4�X����mw3�:S ����;i�a�3?w���f+�X�!�X�3_l�Q�L�y�E�qw��`|�6�G�1��HA�$��e���lu�y�4�y�Y9�N��� ���V�P�"j�3�~ń�X
6`Z_J�m���گ���F�z��w%�ي	�̿�������=EG%i�{u�o�&_���nl��]�I7j9V>�n�m8,��@��Fd[���Z\$�G��&/��	q�3=��!^�K��\��ur�w�N��y�'�Om*;K�� l�w]b���\�j*4`ޭ ����9�˝���!�b֋&/���`�0�R����C���G,� �p��p�i��YԞa�o��;i4c��,��{�����bp-X�o��R���t�^�S.ZE$bYuۅgc�z��ݞ�zks��Ue�܀�:��#O���4P�o, ���_����x�M[]�w��c(�ݛe�o���Bo����'�������p[��yA}�T��f�9X�`1����J�6=�D9�B���E-�:-�$���Y�������j� �j%���RyZǣ+Z���

�B�i�ubƶ&��F$�W�ȕ��N��\�)�yhqE�[��{�)��٠[.U��*��#C�>kEM��h�����4xK�i!�vI�7_way�oV�\��mS�ѫ�eҶ~9h��1� ʴ��;����Z���ɔ*I
��&SL����h^���cǻ�0~���';Y� �V�l/k��@+�ڧ��_�.�%`�	Q��߂���~t�(Q�ʼ�M�j)�2T
B4C����#�d�պ�e{Kn��3B�P�,���>�f��0���s����}t����-��y���ԉ��H��|+Kκ��͖�C�zN���E_��>O@T����rP�+=M�Y�H�[ӄ��Xv��;���R���a�.ġ/��s,��;�\ܛ�[��<{��O�_�ohq��r/�ߩ�.Kt5Z{Ȣ�>6ma�
`j������vf,:�����p�JO������]9zpDyv��fN�;�+r�4U�5�J�_	0g��i+��kx�Ǳ�3[Qu��V$1W8F5Q��t��t�r��?��˫����̥D�u��x�����Q  ��Qb.@��B�2R�=�v�R	$� �*D�9��CN.��VY�˒��oM��aKB��%��#%9�'�����>�(���T�xj+6ՙ�(�Z�c�T���ci�U���uij�0su�����Yꁫ�I�r-H5��$l�pd���.�ν�ʫ�D�\�u�U�1��lU�1�8�;��Y��fa�ޅ�&Q���Oe?$Ǚқݾ�"\TYhq���c�0vv���-�DƭW��5^�l�{HKۄ�Y{�pn�������O6�J����aG
-)�d�*�p�ň�!�pap�!7(DX�uP�HSx*�K��\S��!��2��ס�J͞>7��.���)kY�_�����g�8;z\��q�1�j[��H�zu����T�Bd�S��Gz��4��>�>L'�l��E`䌞�������-�V�5��Y�4$ȔH��$#�0]ܭ��CT��6 ?WӸ+�3��Iz��wL��Y�<������C%1�I����lVc��狚V��\�	CB�!8�������omR)P�́�2�Ƀ����s_Va̚*O���kN�0_,w�v�5a'|~~&A>?����4i~n�pօ{n4���:if���ȭD,�&�I&���S�.�nki�2��^����Sx��t�N �R%�X����E�j���E�_{��nf��#��nѿ�@��r�}�#} !!>�!��PZ ��9�|�����57�ZZ��j��1�ʆpd��=�5�kV�#fFM����Ncmσ�S~1w/��i�x���i�ʝ���ǑPv���6�����[a��G �
�@3���L��a�Y�K��`�"\�q	�l���X�b\[X�y����N�(���W�$"&)�<�ٓ�?��J:��r�vk�Q<­.s^-��hL�cc��HH��oE�1���S�-�!�*����]��[����Lo���k�w���ͦ��p��=��
bV/��ѭ��U��Q�k��U<+/@߆��U�pi��a35=�¨�.�r=�eF�C��o�[���^����D�����!+"2��B�U�v��$���&X��A��TFX�e�5�Begd����3(�3�r	.{**^��gY^��u�S,B��I!�	��{�t"���P�O�at5�Ģ
Bp�1bܭ9?^�p{��z��$���u��A������ζRG�zl�;H�6E�TV_/��	��[�j޹�E�S�--*R�T�t@���f�0��y�Z����_���\�M�/�;M^�ޜ% �R~3ʠ?ʐm��Ss�3p�ϲ�[�&�<Wv�tOB�z���@��RW�$�Oם��LA�/,��p�k:��j���Z�:1���ے�c�Ť��Ǐ�-V�Z��]���>�e_]T�v��]�<�����	�^��:,?�^���*x�MR����A3��F���z�>�ų�{M����@,�N�}���q%b��ם-�.�U�Z�<���sH����(�"�w�Y5 t.�z���?h�Ð�_�o3��c���.1���D�Ќ�ij��K}x4vr ؒ�D��R�	�~M~働ݨ����::�$h�b�Y�$(x$45V9&I����ol��6xF��Jt��*}��l�K�F:����5�&J��s��I�#���̩xd�i����4��I	Sq�d-3����56���"�k��>+y�{W�VrB��� �MB�Z�h�p�	PC�[�����Ԇ��LY'�dG��Q'�ҮMz�Ҧ�4�P �\LB!���W[��Òut /��(��h�um��˛�`�m�&�c6�莅4C�)�6ł4Rp������H�8ɟ���V�P��OQX�L���|M�АHȔC�q'��G�·�3��ʧ��ڄE��@�hNy���|�S�=���A��hT�����}��l}�ڮ��x���Π����9�Oo�Q�[_X;lU<4��;1�]���t���볣L<���V{��,��	��O�x=2b����f�$�c��W={�r�[ё��ߞ�^�����G5����r���]�"4��fu�+�|/vl�q������S+��J�󲵰l����.d׸�fq�4Q>˷��~?�{�b��e7Fb1R�Ϯ5����uoe�]�� c�z�X��^Ǜ��!��Ѣ &�la��g�n,��.�8�+i���慊B+��Fݹ�S���6Z_��u~��'�A��͚O+aUx�H�5�z�����Kw�����w��p&gp��i�y����="<��z5\�=P	��j��f��o��G!��g������C���O�)��c�� f������F{�X�'�k>&�9P�f�(5�6�B����>������6:�{���"牴�rU�7�0���&>&��,��	��V�q�I�4s��h�
'{q�u�;����>����|�����N����Y^�E�-|�B�&4��v��K��mB>ҿ��γ;�&���p"���^�΄�X�:Hޟ\]�5$h�݅c��وz�����%�љ�/�tz� ��5�������m��)�b�^E3I���b:<���������6��E�~)F6�g�$�ka˛�&=��Ĳ�*�hcq���wgOj{�<����Y�u�AE�������/�/�ͅ�qa�sKx�:6�����"�\I�.4�W��5Z���۷�8�(�$���.,A[�O ���Ѽ\d��r���'TX�̲�������ΐ�WOz6��"��.i������A�:�`C�A�������ۍ��E���V^���_ݘ���}���	Tm0zB�s�L7`�ʡ[o��\�J|�[\Ӯ�Z���ɛ�Q/�������P㐂���*6�V�������'}t�V��6�$�/-�y�Ǡ��9�4�x��3��(���>T����\�1���Mf�O޲�k7�5��m��NJ���.��R�C^�X�+'k�O�'�1h�Ij�΂�2.�U��ß����"�l�� J/�k���[E�7�Ugs���KT� �o��:.p�Y4AQ2�*��W��G�t��3P(��ş����BZO��5M}�S:D+x��R9�q葹��͌�n�]oi9� _�D�7(=r�SW|���s���	�<�g��Ź�0�|;}=yvd���G��k_��Ә+�b��C9;�be��8DC���'���bJ�2�3J��õd�.-�>>�|>�C����%��}p��F�Z.�_���ߣ,� ���VU�����>�v�}��ơ,]3˺��I��I�@�'���[�L<R80��4z�>�j8�H�r��a�lo�!L����*#!%�S_������� ��߼��d	B{;�p�Ϝ�Fw�kU��I|��Wd��H�+��o͛�
8?��\9�� |�3�s��Y
�:��(�)�5>���x(�	�cCB���V�>�AMZзn�����|�d|^_���W c�vz_y����jf3����։�L�C���]^^����9�U�_(�Gk7�x��ս;�:��T��꟩�ޤS;��b4�<��Y||�~Χ�ĥ�T�rL��(<��H��8ã�/�#TD�±ޗS�rŢѭ�v#�9AyH��Р�0����&�'N+y]"���M��s� ����aF�]��{&�����c� 5��z��W�|���fD���gZ���Tn��_��DȐK�����5ї�;ԇ���K�"�z�Na��S���d���l�A@zo繛p݁~��u��� ��';����y���=�-̎����^��H�,����+���kg9��I/,�m�,���Ӹ(sv:��䰷evDy��0�A�������z����W�ϡsJ�%�{C�V(�!���;�ó��ĝ^����߼T��E���H�O�*�֚2�����*���5�3��*��P���j�C�ٹb+R\c���1ⶃC�=k,�E����Y\�)~��NL�)5;�,)O��,8�
�EKO�S���w:�H���@�G1��������&AT^��� կ�D`&1��z҆'��m�z���5���og];:��㻙cs��{8��	.�����L�<َ�`�󃋂R%쟛�y�|<��ne�Z����,).R�`�{w��o�~��?���Z>��=t����hiM���+�������f�?�� ��"
����OÂ(�V���>͑p"�b|�G�B�]7D`0�v��S�s���U���_�=Hg�!�R8p��N���#�Z�?^��Oh�Ys	�*&�a��J��]vp��hoSD�!��z9ś��G�F��2�`���o��k�1���VM�%6��M>�O-��0��P}A��3Jպ�oʈ}+��c��Wr��瞨��W�Ê5D���r&�۷�^���%�#	O���MӶ%����;_�OhJ����PN�i}�|�\>(�	E>m��d�qK�*3�Ṗ@��u����'��������3l�D�^��[Un�iY(�ʾ-��"���ug�o������ *R��{q�Z�ՌX�I}���3���OCG6��zQ�\�/�eo�Ҁ��cID�z扝���W[��
#**�sx�MC�wՕs�mږ�<f+++;��,�w)g$`����K��u� CC�U�D XϞr�T�y��=�R>s �<��1c�Eug��d-[��\�����,y�s�:Kz�E���b�K��C;��Q�{�)��Y��.<�x]�fe��Q�!���/M��q�u���6]gOݤp3��OpW�?9z{�N�����J\�>�hԣ�&�<z_�WL���-=_�_E)Ւ��e��06����~��9�O�<�o�˾��� C�F6�����{n�;�o�b&��F��j1�a�]�W��ց�mQ_��*#{�,'���Jn��p�Y����)�U�!D��N[�j�%~��)a�,�k&8`����{vV;x$"��A���,G�`5B�uV��'PU�]����"��b^Hv#Ὦ�B��z��v��Ω�}��\k25}A#�5�d�v�Ka��
Xҭ�\��9���]��C�}�(�LI�d7�ܘ�5�h��t�T(!d����Җ����_z���Q�u�F��H�X
}��8�Ѿ��;��S��q������?t�G^01m�������_ϓ�}x;Vs:�k���0JnHԃ�p{\Wc����6�C�����p�3�K�]���v�l�_�~��鮙�k2��2����]O{������D��O�Z�0+o��[��F�p�nf>��K������7;l��T%.���bO����-G�y����J�oBv�V� +���-;���(��h����S-�ta��.���*���CR��7����+���ўK�g�q�>�E!'��y�kG�?��d�
,�5pk��k=���"��W�]ʜ�{�6�,����3����Yؒ3�aq(�v:<!}2�qW��
<c�p}����\�
�l���Rb_�Nr��)v�_ǲu=�K���!�-@��������!�!�ww�ww��p߻�[�Z�议�:�{�}N����)��b��E�ro��Q����%H�,,(\4��|IRQ>{�N��yD�~m�N��ex�2�ħYy��#l\���o���$�T�,̕�<�h�I�hއW(}}��]�k6�R�OF�5Y���fd����*k�e�h)sg�j86A�x🪰��}D�������9��Ш�@��%Sb��s-�}wQv�	u��j�..a_�9j��(�8�4N�-x��7���P�Rz~�>�g`θ���]c����_jj� A+��u��Ҷ�IZk���x5f��nOBKowJ�N��m u)�~�j��#�F�r���?*��1/�%�0��m�����x#	ք�w�A�;�
ﭘ���x����/E�_�ʎ�\�G��aO#����BJ��Yc{�ٲ��qg��� ��"B��1�Z,�{ <�D�5'���'g�?��������I�7 ٫-���J����~q�j$B�rJs��X8�`ݭ*����jv^�p�L"�d�P����D��?��S���Z��`^^���l�iO�󈡑��q9U�*���{�_�w�?�_�]��kP\��X[z����$����G���0{�ї$(ފ���2y��I��PbO�s���E������ӱ�'M�[��V +�*�$ύ�/�N���T�*1XӚ��u�!p'�B���Oز�) ���Ѿ~���u�՝T���lj��:+n}�Y=YQ��e��$�lU�K�pH��o	f�GJݗ�Yy���2q��6��|�o�Օ��y��v7�����Bk�[���?b�E��/Aܜ�
��<Pr3T�S��Y8Rr�2�m���8�2b���w:�n�;�/b��~��q��&� pu����ajͥ�>�Ƌ�6���n"��+�~�d��HHߍ�f��d��w�6Y����[�8��O��c��X���q���͒��B�[6KY*�V{ΐ��`Q��L4��Su�Qqc_J-Dכ_^9[��&mm,i�F6�I~���:����3DP�B~�X�g)�^7w��+]���i|�ݬ3�i��� �s�����R��P�|~c=~��5�D�EM��.�ȈwC.M�P0#1(ߗXjX�r[�-���+,a�1�?�'�$L,�r���p��x �Bb�����������<B�s6 Ŧ����w�wu�`ů�!�]g����X���z�%!	uW�Ig�<�0�����^*�E �pUd�FOG�ץT����O����U6d[�������'7�̆�22�:�O� C�� ��PC��
����I�ӿ����E���M,_{�	��6�k�RC9�����n�?)��7`}�A�mO����T�W��!'�ˑ����2t���"m\�ݖ.N��T�|O�Xz�8�nO�\N���9
�.e��}��͛Z�`���y=���$�k���|��_��~X�ǻ�dL����OoV1$]��z�����j6�h3���Ξ�˽̑�>���ۨN�ޫ�!F�ySїGi'����B����ć,:k+>5�k�s�Xu_�43ĩ�`��L�H��	�Aa�gd�ylp�j��a]5�u���ѱ=�Y�%�*�e�V\D�d�S�Q� s���-rg׮ė�\D�sz>�}�[�@�A І!�e"K�U�b�L5Q�V�m��W_���.G�� ���� b���i~�i=W��/ ��߃��N��������Օ1�]��c6n���i��� �������dl ʨ��l_j�2ϩ�U�eJUԘ����+�}��I�煛T/���.p�����}Z[m�ċ���>r@���~ʠ��^J���Z;���D��L���B�)�2I��d/B���/�o>��p��@ _͌�Ny��-@V�̅3��ʸ�8��6X���E#C�=�YW�'4���J�f��������{�O�88�w��$�F�Zxi���`����Ѕ���!��SVˉO'�&0�G�kUd_HH�yC
�+AN��߉`�)��qm���?��k=5ɺ���;��	~��
|����~��n�'����s�U��c�q;�{�;C��=^�k[�Is ��P�������~D�)',����;�����)�Y>(����t�@p@o�n"�N�T(X|^��L�΄�tޤ��@���掶��C���q�����&y�P�ki�n}�3(�D�ZI�5�q"r��X�Pp(�Y�ZD����0	���t�E(V�r�ݦ����cZB�����[�e�%>~4b̄�O@ұ�}%�W�Sڼ�/w�����0s��}��!�_��i#�C^1ܽ �_]�;���bwM�z0z<���r G�'�?Zm�h��/]�S|ҳMK8-1Z�l���A���.,�-��榬�f���qX>B�Q����[�u5|p<"�����Tz|W"�7��~+_�|�1B��=�7dzj���ۧpgX�ᶳ�k�qK�{m���ө���=���?�إ3:��IK�ɔ"�	��T��v��qι�PFG���ۍ�<����V�u��$fJ�o�M�s㭝����h�n�J�rO�Η�s���zF�l�+��o@rK�6L�������څ���4@{�]���"���-���� �Hn&V�fNA=���c�_�]�6�z�_y���=���]]���w�]�F������VLX	6�P�9�{�8?t"$�Q����|�ƐJM�Q��E��:��M�a����������:�����y^eR���X� ݎ�pM֕�g��
OO+^%fI��X�/N�{t��
�gA�X9=���sn�F�$%V�v�,P'oVof�#�7S�|�W����Cu69I-qX�0��Ƨ�^���.�8Զno��u��#u��Kf����^q=�G ��%6��'R���/��.p��7h��L׼@�R+��|��r`瓺i��È�^��	�z�gM,�ݠR�Ul�x87,�a���tD��t.F�p��{�<h/9��C�J~���/M3�Zf-���a��ٰJ�"��F��/U�p��}��!X�
3�b���O/Tv}�lx4���n)�F+ȣd��v7�_t~7�;��x��|��Z�y6�V�/	��X&nh#�����'@+u�@��	۾��L�d��Z�����``��M��Y6�|V-�T���H��	މ�6l{����i�i��wn�|��s���]ZH�����\pwG$_���+m����T����2h��]�x��(�h�}�l��"(�pݴ��<����歭IK� ��!�H�dh���1Tĝ�l���V��'�K���{u�w�Ԕ������kX�=�ݛ0��TLn�Z%hj$�e�$j|(�Qo��ΰ����[�-%������l ��͆�_F�{�ԍ8#awi����Q�._Cz�JԬ-j��B��j<.ܩq�0��41q���vҭU�������A(Q첂^��f�x�~~$�j
=�t�(ߞ�����2�=>(������024�?�����E��Jh&�4鄷W�Tpk�4>	?�Q�%!1bӐ[X�̒��\�����h�����b�)�7�F�2��G�g=��Z�Zn0
�-}Տ��4y_���|[0Y�2�n�#V��]�I�R�h'#=�))T+��/�k=V9[)�B���C�l�3���� ������Ǧ<Ww�(��~�vT�o���-K2ԫPŋ��fF�f�b��t��-��"�_L��zd�	����0�`���xl^)��p�h1�q	!;�t\�I���*��3Nǋ�oԩ��>X �l�Yi���ֈV��r���y����!�3�3�L���G��]K�&�7UUDt���ܜ�II�<�����܃�o�n�����$�������J=k�͖����b� l�킰'��(׃���VȄ��7�?�D��,�m6��{th!���86!�@��{�y�^F_�j��ʵ�y�X���D�\���H@�Vx�x,J��	��J:0I��˜��>^���r!��[��U�:kV���Zzr��C�s���p��ms�]~�������{	�7��Rg��v����[T�O	N�\WF�G�q)��/��dHq�J���(�h�[*2�TjM*�%���>��%Ө�
+7��p���\Ez��X�F*���`��Ҧ��ꆹ�$ݥ�4���lV/�Ɇ��n_砝N�x�WW>�ͽ�D�r�Cu�o�;������O�]L�C	�`�M ��18k�v��tt�m��ͅr
ʀ����
X������I>�~ݤ|���m:�u��ԉ͘���V�3���`�H��gi,�~����'Zāk�+�en�y�F(~�'���3��|E��;_�,>Ƣ�͗��Y��k^$?u�I��ok�F�Qي�|�b��0��*'��
E���߯���m���Wn��t~��k�����	�n��;�@ܣ0��x�$�i��� ,ߡ��5�T�1cX
oc/�[�I�?��d�q<��os^�}O:%R�����Y�/HĶ&h�C��Ns J�x;,m�Ӭ��w����j�F�[�WG�*�v<_���>'>���m=]�dGJ�.}��3�%��k����m��MQzD&�����@Ϣ�S���n���\��R����`?G����)�������pr(�j���_s��wHP�r�W����~Xt*$	U�5�yuB�䤢�J�o�Q�7^
��jkf�ssfР"���z�{���/.� �/'�*z)�3 ����e�T;��tz�˭~�"uK&�Q�j�7P��t݃��'�B�������4Cz>ܸA�P2�|R��Fx4.�?�*�LW�[Az�	�fJ5�Bs���]<�n�B�:T�W�n'�/q �e�����HW��$���QTQAhY���ÁҮ�n�Ò�4�7m��'zZ;�=%�֣W��tO��HU�e�8�����롪�����6����e�\Bji����j�Qֵ��c�9_9@����i���֔��Ut4���(I|Pv�/�����z`��.��{[+T+	��E����oO���ƹ��T��{o�a���3����rP�Z�o���U��q@-p�;�'*jC�X�	d��n�BF௡]��i�?86�s㡔�H�t
��?����*n�$E�M��O@���bSQ�.���iHܗ:H����i��R�cj�N6���`�z��/�|�
�,�Ӣ�L`!lT�q�r�d��s�5��t}wJ���Ы���ɥ����$����i�_��Y���-�Ii����Tq!^	j���wP�Y�Km~�1ӥ-�{�5���w8�(�6��侖U$�x�6ԗ�'d;fxAn�1�]�h$���a�����_!�3���
Z�8�nO��qr#����d	�u"s�OM�����a��7
责��P��EY��Z�sd�u��`3��I}-0��4������|)�(z��y�D�@>eq�2����R{IIɺS��{���D��߿?�s�-��9��aw9T761��
��M�@�7O/��D�F�v#ᭋ��z.z��!��[�Gb:<��Z;Vc�~]_��D J˲��[���4�����}�{�'�����/|��nQ��+�s��3�zm�.d�	de{"�{PR��Gy9���(͕H՚��K�WM�mw35��ꁢ~��\p�O��u> �[�3�Z�^�蕃�)��^��M�N� �ފz�Р��rg���I{��됁�
"/S�Vnϧ3B���sw���[�~��'t�0,��OPOnV*.)�k6r଎g_@-:��N���ee���u�7	t��1QPP��㓃�C.67	i�ݍG[aiiа��7���"�CI�-��럠��d��g�1��ec�ૅ'���jAA�uggN(��Ό�u��W~�Oqq�KO�������H��Ә!��77�ƫ����h.�u�e�*���u_R�u�ܿ<�!���aXܯ�VhR�,zW��z��m<!Cb��ú;Y]]�ڝY
��>Q�#����c���5����c3�{*3%�Xʏَ���C�ږ	�N#W�g	�P�e'5΂ţM���9��6Vɪ��܁�qh�;	�׸"8���Q�_�C���^�U�1�ϝ�>�b�Aɚ��qJH�!�7[�ړ3�P����r~a�����Jt�B0�qF�*�*dC���x*A���@p>���/FWK-��7�y9Ý�ȵ�l유��<޷��^��}`d��k3��L��G��h�
�\�%#���d!� �de-!,F�|f�����	�xZ�V
ʊA�����lGP�y�M �aM�J@S`��l�I� �S���Q��P�<�H��ED;nob@R���]��tyvv�|��8m}�����qkbya33H���-����iX���D�V\�pӤ��4���= i�\f�&��U]b+6�.�[��E=d�~hg�zbV2�߃�N�����HB����z�.���(>Lf���0�5L���M K^�O"7xV�n�`��/�� � ��zX\�Q*ZwbX��Khx� �@��u�;_����0`Ѥ�5˸DA� ��b�Q��ّ��@㩇>$��
܄Znr����C![�h킽q��6�n|�E��	����?� iyyͲ$c�ެ�}ů_����9R�����Ao~֡�`�4b�*�@R���Ymxf�q%//!IA�֓n���3�4�9a�*鐇'�O��wU!��f���?�^���\��-h�����K@HǕ(����!A0�󇃘X
�mE�#z�ڬ] ��A܍��"�����h����w���| ���g�d���T�Ǘ��<�.o���֘�~V�uח�H��Y}���p?hb*TM���l���M�,0�U�J�*i&�c����J%З���ʡI>e�Jr�i�i�D�^�յ���y�G@��������ԘI��V��ݗ�=0�Ë|�и����7[[���WJ��2qn!��D���#ڃ��P�(E6ֲ�dzf_<>���*\u��~�]I�d:Ne�5T/��u��Ǵ#�����'���6���˰��w�Nx�"�Z�M����p�'Z��>�='��^��
	�K{A�&ZZ����r)��o�M�������텳�4E?N��4#�����C���#_~%-- A����H.\��1W�A�SK@az�� \	0�Q0&I��\KrH�.�h�Ń���\�$������Hފ�Kȟ���;�tI�
ҳ[�_�5�4�mP m����ec��V�燿�����G��L?u!Y*uͶ� K�����M�]T�e�\LcM�]뺣���ބl�~)��e���\�w�3੅�d�:���`su�sP��	x�.?�'k���da<MD)n:���[��:|� n߱N��=��}r/y��]��{��I�z6��N��B��nV&{Kj��J�n�[�t��m�`4�K������MK;��#��m90�b��2=M���<W����l�tmh��3{��6��k]��==���>�O�
�P���y��Hg����4��fӡ)@EݧC�Zڵ���S�z��Wݷy����k�ĲE��C ;�6M�����	J?v�z���1_��=�t?�#�_���r}��c�[(�&1M��a�D�{�YMB`Y����rj�Y�d\�D��8�g��d� �	8B$V�&Ā��Zu0��A?��7�-#�P�ׇQՆ7�0,jY��������}�Rrrh�.Jm����k�!����t��H
�A���wPjD��u�7V�u.�sٽ�x�oJ�Vk��X��6s#a�?��rp�]��N��Ծ���3�f0G6R�q&s��^�;���IX�x�c�5 �ҕjv���V���N1tF��M䣸��*:����������#6|Е@�jzï�}�V�5�]M�6��5�?¾.6�;�y{�/H8�FN/����O9�Վ��Y���f�����>5;�B��^�S�-C���]\||w��/���z��_��� v�G�Ḹ��+����������t�̓��3�0�$r�B_�/uJ~�dKT/�Y�̋�|�L�M,~�	1��K<v�R���W-ɞ%6>�fθ�m�n{'�ˢd���=�����ϐ�X*�-����~ٷ���OϺ�8r�c�8�Gٯ�ct_K�a\�F_n�5i9�2�Z�gYQ
���M�4x�����X ��^h9�O��D�HYJJ���iW���]��KIw�gD\�)\A�1����+-��)��S�y�H�ǚ�f���=��]�ǯ�f{nA#�o��c��F�y�\b%rQec��<���@IO��yݷJ�ƚT�<	_����u%�+uh�<	��ҎL���=�'CU����c.�5y�}n{g����lo; �Ђ1}mӿ��x�V�EU�%VC�g���d�� ��I����is�鹵p�讘�����h,���fy�Cˢ�X�n���+m,�2!���8҇���aS1�R�����Ǖ:x�c�_�Ҙ,�X��X��λM �A�z:�j.��]Cm�֍��4^��2�1^QW�n�X��q��<K�T�ë�Do�d=��zƓª����E�dO5�E�%Jx�c�����m n�쒍/7O>�n�@f�%���SNN.5f֝G�CY�y�)nr�$���t��Q[[��L[<m�^6�,�7cq:r*�Y�)�H�:���ҽ�X����c����ҩ`
蕲[x��ڧ���z�{�@�+勠3/�8����	��LgX��Ӂ����0��7MAf���bYx����P��	+�h�%��\*�x��*�9�H�9��8(�f+�7w"0]�0/��>*�����4em���V��S3���/�~�X���AWe����P�ϡ8�cl,�Q����MC�5��ޗf�#c�NFg���f'��=;�8��nH`(��7iiT��o�[���b��]������@d����<NR��g��޺�,�"�L0!!�";��A��8����ts�5���4 IF�%:uĿ�h*��b151�Թ�����^!��o��A p7���e �S�q���zʼ̄w}224����^{�"��%wv�#5ԣ�+�=�U�f�!09��ʹqD�����Yv��W�pEPW��ȃ����@�3��n~߸FK���¾�e��2V�夠� S�a�DT{{{)iiQCC*&u$H"'�^f8.���ϓR:���B�� *�Ɲ���EǒZ�C_szg�D������u��S�5�@U����A7r��*�O�k�':�k3{ ��͓�5�����:�(���|��9,:�֕��"���C��Z�6�����̷��5���mQkk떛��S��׷8gF,}��C�ڗ�[	Fcm��C6�畈�c�6�׬<0�~�F�S��l��;�d����T���>x pK�5M�-�������u2#OII�RP8Q^������O>+��|�h��x����]@Zb3{pŖ"KJ��$ďM�d���V���1Ű���V����兪_���.[� {�^�NG�y�Ւ҃�������l��0*���۸��]L³���H��3�>j���k�9إɼ��v�N�ܱ�'�B���t���nro��QFZ���M|��*A��܂e��t�c�k�*���߫?���Wx��,fQ�$p�����%{<r"�����U��h��fh����P���ҕw�m{3��<��1n���ݢ�_��5=d
����6� ~��m;0���I�eφ)��!��"��̈(���b��O����~����	 ��1��E�p�U^�e�\��o0��r옜˜�Nw !aPhE���A�СZ$z�d�Ӯ�~�}�j��͓��>F�Ǉ)e��>���Sd~��fWBU����k�E0%�ꕔ�Ⱥ{�t���	��
��AI����Wp!��R��`�x�'e=���Q���D�O%�.�`�����o��a�V觡�sX�3����b�<�#
c�0��~F��!<��g	�U�(bD<��@qd�D�Eʶ߂l�mE�7�F��*G���gZ���\2�����i�.��t�ǐm4�wv��w>��SK �W9�@>�5�r��^�<�ۊ��mW�����dK��0,Nc�_����nݡ��N:��6����s��9�X>/��
�)Y��1=����@1;K�h�!��w���H��e�����+�@�����HH�.���"۟X���h�A������(�|��@X%n�R�ӹ�H,���:�_  ǎ��\]�r�{�#ztt�f&���?�[qxI�i���FSn��ٍF���g^�\
+��s�Dҏ	L%��~BN�'��hz���BsGJ��q�Ax��j_6�E�[�`"my�^�ki��j��j}8�B�;��� ��HY1���hl���.g���(7e}������C���	�F���	R$@����p�s'�(��42�0T�Ha]VI�]�Ih�u��1��7�ͭ>u{��~�B���g|	�`�������>QB�s�R�m��L�����E'�|�p٦ث�h�FfoG:�ݻ��;��k�]�{8�J�cߺ�<;S(���~kZ���Ï,��G>+?���V�K�_*��w�h��~ե&���{��޷be9�
�I-ض3��w�oZ:�w�wz�����7�;O�,z�Toc
/���
���#^c<�A>q�zT�w�Dr�����)��-z�<�$�D�����?�Ћ����i����S:G�4��H��Y��t
ӌI�� ����8D*�۔�.Ҁ����Cf%n$��3�I�p��QAAE����:	�a��j#�R���K3�i2���9��~G=��]��^�[�Y���,dAV��-�X�κ��(��$�����K�o"=�n��u�^�4�X]F|c�p7hj'���"��VBo>���s_��W�p�#�����6�������O��<O���׬�p����ko���\�ڗ���Qq����=�hv������Y*��
��~5�S�qlc���׷���x9f7��!��2����0���ry��0`DRH�Pke��{�I�mC'��9N�&������;��w�T�	�-����O�hkHy��4�wz+hd~( r |��l�2R�ିr�'#��V�^W��]X�77���5\\^������D{�[��u
��dh}�+E�h���l�v�m*\z�+��i�!���.��[��{�.�}C��L�/�#v��%>D�3,ߵ嶌�?�S/�؍��n�Rھ7S	{o��&H�,/,1L9_�=!���#Z&S_S��į�j��uMG�x�����S[F=���b�`���A%O-yE��aĴf���.r롼��� ѫc}b���%OT�S�|����$x�uL�tH�b.�r4Đ�À�q�8zCNNۤ������d�Ц}w�+Ӯ�<�����.[��A3??w<�{��ܬ	�HF��,D�L�ϟ�H0�Yn5.����@���W����@�����IN�А,:������@�߿���>����[����6ˈS��dS��B�6E��?�~��7B��� q��=D�4�U�Sq ---���hVmk5�)d�ܱnL�+_���;�;�j:��w\p�+�N�w9֜n�F����L��S?{L���7[�fv����?�pD0}�iD@
҂�*�g>�ʰť��B�TK8��SdÃ���1����|�`��⢮Q�1II�e��w��Χ��~'666���̗�iO\I�Ȁ��a�q����+(+Kz>��,�|�� G����t[�H�Q��f�@�?ZXX|�&�Ņ(�7Ӂ�~�'N�?���HL4�{p��r���1��_r��6"N _3�a��\\�8N�h�����֜X�t������1qq8ϱq��P�+$$D�@�'=$^�
���#!�#�kfT�w�I_�-��{{�~���>�g��al@�[�|o���~Sq���e$�GB���k��}�z���$�o�-���_�c̑�5^�"!k��(�H	b������ۘ����<�z�XHBV6�T�C�bb�
�?'0�Mkxs*t�_/ggg�P�%��ı��	8y�m
�����Qz퐏�N�P����E�}3���=���#����38��7����g��B�F��V�w��hk�2�1�5�TE$Kb%��)1�|�T̤�F�K�/\Fk2�� �lF'�^����B~D����"*���O�f�}غ@v�!�DQ�Y�#�e�;��_ӻ&�٪�nް:BfS$;�r`1w�9�B'�RωB�%;����8Ce���Smr�
ꍷLyKWz�U���ů�@�4�i��R�dj+�wH\��;3��#�&����l��?�PIT��~���n?/pzN�y�M=8'B�?u��!���![i�-Pa����t�ko�%�z��P��sp7�Ġ%�a9qv�&��^8������*���<�~�nu2��\M@������|8�<�躎5*������[ ���X��[��ׂ����])�l��c�k�1`�l!腳����\�V�|ѿ_��yǃ������t���۽Qe�@���4# �B]�W�u5�kd�Mi�l�v&U۸7��[�Qͱ�����ӳБA��/�0�,��E��t��[�����^`�q	&W.�$X`m�}j-\{v��&y$@%�4s���-(L��B^s)��X�E
�^35M���X⨝��[؁ۯ���s̐�4��&];���� �Ƣmɸ����ӟ׬��6����dmG*u>e�T{(����}Ū�ZR��柘殢/��R �m�]�����00���̾�H�r���^�o�>�վ�.e��]��/y�����y-��D�-�����Zi�Tf��(��0��Vg.MFa$#�b�]\���Gv�P��u]���T��[��+(�K��A[��B���]�V� qX��(���nkx��uo��RN��Vc�ؓ���/�v�{��_���<ڂ5�����$2i(ܪ�%i��Z���z��������L�A�k����5�k���AP��5΃��?ɲ�ɑ���Be�n�x�h�Q��:߲g3׉���II���ێ�����L�{K1�SX��	��{�r�H]�R�^���m:
d?��.����*��a�<��p��y1��F���/�B�wH�����H+ƪV�NJk󖡯+� @�_���a��s�ˎ;��O�������:A���b���BWP��fk�q�B&�Z���NY���3dy&�gI�f���T}�OFܽ˸��8�<�z�d�~�Y�RT.&�����j�$�Nv+\3@F��韯3���gų�2����8�ti(H�����u��rQ�u��b1.��3�7~�8p�q+�&�cEJEP�%Wz����[���o$;��{S��T����^)�ʏ��.����� l���8i���hJ�d�_�H~a7Y�B������}B�Q$�u��#�w�g�D0�\�����V��T�
����jN�{z�Z@d�m�dX��s�t��Ί�*+���aY����I�Y�J���L��%�FT��;XO|c�ϲL�:걕�� �a[Yȴ/������&M������(+�̆��Ð�����������#��gtl�����)� ��X�%C
U�umd\�rIK�"��R�K<Qb��T�"a�)�񇮦\���,��z�'���4s7��I��4�V��+��܅2RUKKU���:a:�@��"�h��ɑΏ�b�d}��v�K����R-��p}����ʊI��We�H	��Y�m�iE�C��g��]�oJ��� �Q�?7����񽵓r�PX�aH�t�h�1�ɴ�DH�o��0��㾠��f��EX���j��<�~�}S7gs}��ٙ�8���o���n.E�#T3�n���-Op�ߛ�g�$�7�p��\�F����DJ
L��;G��f���`��>%>�#'pgys/m���s+c߻�{*���ysN�l����XMGī;��.މ����t��Y�@ǽA9��Iۃ�l"��l�����1�}T��� �O��P�~塨��r��>zA�x��&_�f�>==mm;��.�a�lټ�;�8~�")~KUw�\̝�}JI�I�z���5�G��<�^�5i�~�@�3�����W�Z����೵�Xq2l�4�i9���?ؾ�x=��?Y�s����w���33�PWA ���s���ы�T����Mf<���7���z�����-�h2�Aߎ�.$��6�;�B�V[�|���˅$B�β.�`ôZ{��r�@-�X��߰ ��:�#J_��L��'�떨�v�C!��6��A&�%�������9�H�)w��8����@��5 h�$��ug���TУ|%Z���gw$J 3���k���<+ck�+��Q*�M�֒�?0GJOm���
�0����ĭ�o�jo
���<���G��|wSW&U�82�j;��b�	��������^Ū��RB�Ҳ�*yq���$��X�"3� �l6��45Z�`^n�:�d�B�Z�o>�{_bC�8��=��]F�R��2�ݫ�0ǲFuO�����r���u?� �i6=����v������:��hya�P��*D&�^N*�I�b3C�����3����E��хï�s�m=>7H�[�/U�:X^fc�Y�ZMH�=���w��/���c�������9�,6Anj+7�r~~ՈC8�<D�/�E�A��m����#,�?����?�.�gCC�u�IٜjP��	�(E�.
b.����B���'Y�'����rV[7e��L ��6�ݪ]�	��C�k��J:���B��Ԭ�&{�u��+���K����|!�!pn{�h�����Bb?��)���(<�d��t���>���9�w	��lI. J�_���֞���j6������0�@�cIq�8�N��"���&o��y@�JD\��P�@�}�Y����B+;Q_�w}#�LJJA@w�P��v�������,h�v�����9���mgds�
$���=PG�,s�`�ͅ�����������������?��}��`Nt��d:J/LVa���{$1V���0�!�� :!� ǐ8�K[�Sc� ����{ ��լ�Jf�5��7G �c�� ��|��8��$@���/=fl��c����D�����4�/4`���s
�!; m�%��=Q�+�Jf�%�?5�5�/K숮�'�����- ��q���L���v��1��E�B�9iS��)	fS�&/i��U-,��Cˬ�{�'f(�����l�$�I@lxW�d�R�	�4)A�<��?��|�0���@+�4�l<-�R�s=�śN�<�H�Ӻ�����@�an����5�L��L��z�^��z𔅌��BXPQ$�ͨ5i����B{r˥��,�˗��p��l_�0�8׿�1��DHAA\�5�g�������N�|bK��T�/�7��-k��x5,D TX��W�w>�2��D����9��˸��C �X��	�����|G�b��� ��-�&Ե��6����BMvQ׎!�wM�X��tl������^�!G�++>�l�Tr�5�;��}哜��ա��d�+s��pV�?��Q�q�d}�ԥ��9��ͩ�����ͮ�!���O����MF�t�7��q��L�����XR�C�_��);���q�����S��z=�TMtS*u�$��6��{�E{{�j�qƊO��ĲvxZ/yZ���mG��]#Q�}�����<�L��C�8_w���_���I�Z<�[�o���	�&gcZT9x��lBd	�B)S�>�}�~9g!�YŤԍ�]�$������ܚY�t.X|1Ğ�AnL��d�yFw�Z���,A�\xğ�U�fE��14��?λ&�����n3�W%)��=������NL���@��xi��u��df4�)�f��Y��F�ھ�:O�i�|��d��ߋ\i,�������������TA��	,���o�w�$��K�s�_#Su�#��	��~v�E�%g�3�2�]���g#J�@ ?
���.r�		,Z&恊��^v���M2���O���8C�D�xt��<���,���~W{8빗����z`R)����*Ի{�5W��M�cS������]$��$?�h U���AQ��7��~� Q�}����S<:%��3�_�׻FC��Fm�(J�U��(j��Olۙ���#�}U# qQf��C������.)�Kj�|v��b��h�R����P���քw��+�
�A?�r��o�KW�\��o�N^��t:Q�"r�0�dU�]�^jb>}5z�m"gd[R�
΄�ڷ��f<G|5A�@&�/�hA�0B'D���;�v�-[@M�7�j�L���֟��?�bʃ`o�
�eFC���͙7P���s�i�8�t�txf�ثZ1w��<��U8�Un�!����+��ɥ�8n<��g����_�ѿaUn��H,�A�E�U0��̇�c��}���� �]�ڑo��yR�K���'X�am�Ye��u��dI=�,����<���pk��g8���.'e�"[9P�_Wշ��n��*W:�@J�.����s DJJAR�!�[b�nf��w�{w�{�ޟs�Z��Zk�7Hu��Hd��p4Q ɝ�2��:rl��~zh��{�+
�HP�k�$�j�� a}�������@n
y|��B�/o$�؃�!
C��Z$��|���T7燯w�j0Ù*'���C:M@���Y���(ř�fXgq�T���]шߟ֣�-/����G�xh��^J?R ճ����0=봎�uVF�2hZ ��i���|�����_N�|���"�VS0��^���іx����3�����li�*�I����+!�ny�Q;�g%=p��^D
����u�N�z �J��{��g�$c�\s�ȾBb$dŭ��i����&��W���)R�E�Ę��`Xx��~3�Mk�3���1����ꐙ�%К��*b��ڙ�qG�ڡQF��� ��u�yX��\�6�����2��P,�9V�u����P�0�qX_�h�`,*�u(�c\EA�+D�HF�6yy�>Yr�7�X��A=S��´`-l�OhY$�3�����e�L+-�'�/}2?���������aܘ`�8��W��X���B�KcU���k��Fb����y=�;&�,~�r69�Ñ��Ac�m�/�^��eX��y�$�b���	
�^' ]�ğO��Z�x�Q��-�Db�b��e5��.�ÝA����Iq+0̾����}�Ǩ����������F�GxM��WȨ�F��p>_(�k���l�{nF����/��u �.@��������.��q�pX��&�;�"��rq�D9���\��s�4� ,g��.M[�8)kV�(�~�cuR��!v׊rH���	w5V�l{��	�yI^
2�o��%����� ��o��a���LG��d��1��}s���5-Q�a�.���������DD���6�V'���g2�*�+���1���Z�)6���������Ua�w��9p�{�Xm�sK��q��K�����m�j0Z!2xNzR4� c���==z��m��9�"_��d,1��H6k��
�|�i~����� �?��g�Mi	=%��B% �ET���ǖ�@4�Ϛ���H�NI��hH�Ԗ��8�/�߲��8�y�6//'��T���p���i���޹�W��r���ER���J��:
$Q���
�29䩱 �a��3��<�d{�z�L����q�������E��E,1a��[���Z�Py�Tsق�]�x":PbN��T4�n��������|�6܅���1��K=�PK��6W$-e�E0~��Ŷ�?��݈N�� g:�W ���3�n��H	��8M	�h��o�7׎Z0�'�a������0�cאG.� ⯏Q�6 ��'�*�N���q���:����:�x�y ���a��������L�T��+�b�
�������1�)�ԬE��ܜ?x���Y�ց(����!�`�ƣ������1$B;��oA��a����@^f���!�p%.�|I��OC-�1@A�~q."c�&!�ꍰ���at|7�;��]ͱ����wWϏRG�#W)uX�ߛ�@~�낒wP�!�����u���Tlg�b�	�* T�F7���seW�_eV���n϶Zl�ȭ�K��s�\4p�7Ju��hF׳(����>�Ξ_�;��j�.G���]Պ��/�8RD;X6�;�}s\�#��t�/5|���U�Ҏ�=��?��(H�b�|��FB�f����E)�X\!`�+�;�������ӂ�ƚ��dh�Hp�x��M0x+(���kőb�:�}�S�ac�V�/0C?o�Ҹ8A�N��]����p���]ɼ���_��}"/��"�!m�sY^��eSZ�;�Y�y��}r*�~��%l��X+��
}������߾/#��D\/��P����d�)�4-�}�pM�����d6����MI�B�P�;�$�kfc	�7���IRA���!�f��zZm������d�-�n��9�P���y�MR��KTO�]�����d',�+U�WJ�W �)c1�(W΢@4 ���?�7׉�Bv\řu_���%5ta'�fϚ;�N����E�ڿ\|��n�K?w�%�?_ ��GCKy�n�H?O�5�����>i�^e��))���W��wa
R����k��{���g�u��)��t}~����^NNZ���3����Ye\�ާ��HL|v�i����b�0GrZ�)4�.��0q�_�dbP��`��ԇi����'�R>�n��\E}�����_��Gz:�-;�3�g��3[�#70�7Rp"��a�
U����OiM��}Gk���l{|-�����l��!'~�
�7�ӉRc3Ơ/�K�:K�ˌ�8+I4�o�<���dq�r-D>Z�d,1�%���";ˠ�B�I�fֹ��|1�1�S�Ob�C�G�ȴ�>d�R�#��h�f|��*!6��~BR�f��9c�=/ܹ���Z�mu�VW˜G:C��dUc���9N=ٕ�	](��"�=�V�_����6E��M��RiN�=�i��W�G{�����q�;3
G�]W;�	���ץ$�fw@�z(M`]�o9I��L�z���}�>�e�f�p��&�^�����J��VT�2�F�h}�i����������[yy֐I�{t�oSh�=i0�#k��z|b��
����~��N0s�uG�^�`��]rz.!u������#mc+��q��{n+�܂.�m���4u}k%ƫ�1֟#Δ�.�����������A2�y��'��-#U��(�� C1���k�޿Q�1{��'���:�u*و���%5(*]��S h:��\p�Ss��Q�C���敊0�MUYB2�����wa~g4��H���,1Ѻ�`/ڒ���`-�*\��["�Q&�zH�W�[Q�7q���u�-20�� �pY����=F���"�������)ߖ��mƋ��㝙�,c8i�;*icJ���B���!�����L?�g<�>yM�hpO%��|�H��.������!\{v��ߜH����I:i�\���� :n7��η���}��-�o���J�"�o�������	8:�$��"G5�NU�{�3Ŗ�c�%���	���ˌ�і�& e75����G;�l:����͖E��#�{�sş��鱯���'?6��/&B���;l�h�p*�u��ȵ�58����^�	Z��D�2���	fؖ����#�0����Z�Ry!{�b�g$��8Ǒ�N>��oZ\�0R��������R�R�W��O}�,n�ιZvP�u0�:�����͡pZ���5�[���	3�t�(�yA����>@j\�e���1Ե��wR�U5u�����b|3^����I5Zd����Cl�o$n�0^s:��?������[�l��LU�T;GM�F�چ��>���Ъ��i;�N����$[^sU��a�	��O�P?vmzʝ�{�C'�rbc���U�E�����^��O�ɷ���\~�]N�O���?+:���|�f��]��[q�q�� ��*rk�͆���R��������d0��~?�̇^��{-z*f���gq;��"�ތ�K��.)ߢ<�� ȠknS)��jT�/l����F��/��'�����u��
2���ƥ���T'ߌ��š�bck��~F,�k4a��\��6?�\qO>~Y>�'}T%F����v�޻8�p������>ȚOc��k��(��}�7��]	]��˶ss����<��d���\�r6"�?��Q��3�26�wX�(=�G�I����������Qݏ*�{��̉Z{\��؄��k�`,��\�@\[H�
�xˇ���������0��Kx۶<�������w���T���w�%(?�}��,d����8݅��N�ߺ�F�fTPZ!}�D�z�dv���zw����HP	}I}�2���C�/�r6���M _������Ր�SxNa��k�Q	�����M�u ����h�b.����TUyzd��ӝc�Fa=pk�WU�|�(�G a��]���xx*)r��N�Ii�Cy��޼/�ܵZt�A�-�S�O1؝���^6"oL�}^^1��O�0�q�c��HX�a�����6"�A���K��:.���Gq����g+ˌS�﷞�X`�"B!Xtv���^��5T����4r<M�$����`����k/瞊��)k&���^e��U;Qפ��ne_*�_��+�hY=:�0<���	z�5����W+�(T����#�_�g�>�zi�uj��B�fE��x�Ó��P@�b��?�����.���*"�0�S�bu۷W���7�i���3
W��������aE�R���`0�_Qz��<�Z�)(���o]�4�ƍ!(�z���qJ��:J�,��ҽ���Þ}��Im	
�y_���i��lG�}���{�q�v(���h��}���8��-N�#�ށr;`�^)m1��
�˶�����[w�;��� ����W� �J/�����PK   $d�Xx^��6� _� /   images/3c85acdc-f066-473a-bd4c-bbee71bd49cd.png�e[U�7�	%AJ$EZZ锖��t�tw��t*H� ��i��nx��?�|����.V�9���k,��*Haac�`0,�7��0�vo�>�I��	9�����{}#=_-�?|�,��bg��f������bak�dlh�����,uG�{�QuOۚqsW����~�{��SG��A#��)��C"�9��-���LY�YY%�o4��k05^�4աs��2i�=K61x��������S��<=�����*�����f��fz��%����#�m�A�����{���=���(@��#L��{|��E�]��4[���0����9������C[J�P�>����O�i�<~��@��X�	%%�[�{777����		�S�b���9_f:��/lMTt����S���Ow� �BQ$ܒoޠ�������EECC�̯�q&���y?j)���^�Sk�����x�?���i����N��#�5[�g�`�s��Z��BC��P�<W�����fFF>L�s������|����0߂D�s7M����b��9f�*�
Ӿ��[��X�����VR��e�e�]�Y�$9Z��3DVֳvs�n3.O������Z�9�d��ikC9o��č���nO~�MdU�e�[=8%�+����)8i����2����	aĽ���7o޴4�\�UUU��?{�3d.��}��ܠ!!a��L}�l"KhDDaUP� �S�{����hU�3�׻~�d�P��\����L�/�ʕ}2�:e3J�Q�����x\�����z�� �E��}ϙb���X�l>pm��Ivv6�?�������l�Sn��8*)?�]�%���H'Fl������#���B(@��f(=8iׄ^+�O{�6�_�w9��VB��]54���g��.��d``Шwe沙���~q)t�F��`��(���g���ѽz5R����?����,{�KX�[O�u��!^n�	�3�Z��C"6���951����>#33VAA��~o�+��y�݉^��j��
TЎ7FŮ/��~X�}���b���w��?>�Y8�^Q�?��o8���x�la��Ak�MB����/b!�n��ܕ�,+���x<�����).M�:����8m�ɣ� �p��S�{���\���顡�!:6v�v�\4��ƴ�7l�r��x�W�F�� ����PfR���(�;�K���͐���M_?SSڏ?p�ƥ�E��<�l�|~�җ�9������%ayy9���V0�
ߖ.
?�P��׻%���K%��+���|p�_ϧ722��ʸ'�s19R1�eee�5�:��pFq))*pM�O=�:�5��/�n����*1555�8v�;�1 O��2jJ,����\Ɨ'��|�����S8��Yt��3�vD�]�K6�>*ߍL���a�]I...�mUd�\��71mMV>�w�j9ٞ���YM�ZZ��kkk�:����t�x���q�Wx�jE-xa�O*�<�i������ٶ���͑��l쪚h[�K�o�����H���/�F�a�`	���1��bE�V��m�!a��B�U��<2G�J�ɮ��~�������p ����^�"�]6�f��\"H(�Z�hj�Zfu_�M��m<U;K��ʆ�����UGG����mN�Ѵ{�"�Q��l��o����?��c��c�c����֔A5�Q�W�B����K���ݩY�ƼM[__�hpgo:[|�Q�2����h�=-�������c��1����j��2�ς�R�����ܖ��]�����D
�ri}�6>��R+E�?
�ӧ�_v�C�{�'��ӡ�"��U�X��b=o���"�=��=
Z�iq�~s�o�%����z�-�X�J-f�G�<����U6ڷ���`�p�s��a��{N� @9�;k� ���:]�9�wu-%�������9c�6x8ɥraV�0y{�Y�Q�HSe7��LyC���M��<�S������ Dn<(���D^Cm��z�SQ���dCX8�����������YaQ
tt?UW*�kt�ZY^^H�kj�f�؎��w�/�A��~࣬<|#�u��������8!7�|E�-�$LH}��n�������vԙ6���R��B`qK�F �����̪��m�;�i0�^=��YV%��)�����McG�4J�%pg���Tc�Ï�f�D7��p�����2�­�A �rOu�V�xz�脱6����=�5�z+�}[v3�h[[��c�������u��=������;�gBB� Ylh�6|@�����!H�������j�_g�D�͊�݀�I^NN�8\�P&��F4"<<�Rf�y�9S��n���!�@�4��@f�fis4�t1�'4b�)l�䗹�T=���{��Wh�]8a���ư�Ĵ4�/}����G���=j��_:���kW3�@��O�:��*fDF<aU������rJ�c9�1F~�ލu�?=bO�D?<���Z��j�Gǿ�ᰳ��m�S�+�h���?k�-F�B��nG� ���f<�-A0�	�{{6=�mΣ��߮��� ��f|8l�;���=ӊ�qD8�\�'C6�?SH�3$R�]5���	�^;@�r ���9�"nN��ZH��v� �$qۑs���x��O����KD�2sq�(���({�o-/�����ç=V���F}�J�p4,;���sW���n�ᣟmm�֧���PP�b(X}������M��Tʠ�r�*��OH?\Lو���_\nU��N��+�0���G2;V
0
��L� I���39�2��=�� B��U8z�a4�4Z^���6�6o�mK�������^g�a�z���W�c���;@��TZXK��D��H��A�� �u؝ ��K����2�����6=���x��)�滕�>w$���Lʪ/ �mxsu��č�ad�Ê	�l=��A����2]m�W���~��[I��؈eN[G'R���p{�NJs��P�vF���e���v�䒶]cn%�4!E���7M��А��x'�������n�{@��޷�#y��N�s~�o��� ��;���|?��pGJn��r>)^�g��u��s��>��S����(�S��>��n�]��^�����]��TЁ�d�c�H�2�|t�z��;�p����.@�u�[?|Vz��_O��ݕ����K�ց߿ۃ0����E]��g~w�Q�_�O�e��'H�	(��c�&�dQ�]���fj��ŋ�\�G�F�1��� Q�})�޻��S� N��w3����S�)���h�0H�LN����`f�jDo�***� "��t�GP���lzY؏�щ�=�rI0??��SÃ=g;��G��̠V����; ���	�nu�P�{^H��?���0b�L@����֋4���"7�w{�2���� zz���g�᮴�D����ϧO�+���0K$/�(El�F��
<z���y}V�f��Ͽ�~u~8�U��T�aL�n�b@h�A��u�r�c��`�˔���{`	Ys�c�ddd���	��~��T�'�I!��q,f� vh·G�	� ���*3��M�
 x��x�w��A/+Yan����֖:������{��ƳDP�4�` yRv㔍v�k5*-�� M�HȻ�w�eL���8�
��>!;<22A�/�V� �ǿ�r�|�������)Ґw�)Ԯf�̬��w����d$�iP<M�!W����'��XP��`d���suF>]����=�K����>#��#p�L8Hu�|����α�´?-��i��v�C�WH��������|����}��s�]M���!��sxO�� 8�Y�RP�g{mغ����(
��x�J�e�iW�;����A�((�Sa�0z&�v��F5Sd!ß�G�㊥lҁQY1���@
�4�Vj�{�X�-kգ�m�������Yj	�3�ZVT1P�ͷM�K� �#+;���q�J�$�7�Cl�r)��|�2<���kGJ.����`�0���+$��2����0�����B�R�?:K�������j�x���jP��7�H�{��V]����w�|`\L�$#��ƴh�3� �mPxyD�w���ᐜF�����rjN�zU�W����n�NR�
�MB���❜!Qoo����p�{��pJ�y�)��b�> ���x98���b���w��B9C9���k��/|1����0dX����;�c��׼<�&3���z�\"�T��&j�X��ϊN1� ����{]��(XOUk$�|B;���؜Q�S,�aJ�w+1����]m�ߊ��cƕ쇡
��[�d���c��'��ODC�$s�o���"<;�e�J�l�"#I)su,���I���X&p^�&���S`�Ȫ���
���d�-���4���.�R4����������jՖ�/no.S��DE�f�v)yx4��z�p�� �£��L����;'��,oT�Hqmf�^z������nW���[��?zJ����Ǘ�FC��z-G����WPT��Wʱߙ��J�?���?6,�P ~l��ژ���I�*�4B~e��ރ�%\�Tqp�}	K\R�R���'EHHu�o�f��0F����r夥�b��Z�```$�|�����'�ݞ�w�L�TO�w���ӊ�����½4��rOS�_�3���44�J�J4ak���}`uRM/���a��2
d��bx�5��wSŘ�M}���Ic^��P���MY��/�e*}�/ڂp6m\ >b�cJJBb���f!��^d� �De�^0����;�P�E#���-&���p�%r���K���2�[߾��SR#c��Cf6䄄��z^��K]��~�w׿T�����G�W���.on��ύ��v������Ж%���;��`�|m��b�2F���=C���v&��H�*�� gQ	v�������}Ӂ���5��_��J��Y[[֑$��T߽�p��L����t �777װ4�!�t.�h2��?j��-F�}�����K.���bƳ3�H��	�s�$c����haq�Kr�J1L����K��qx6RR��!������e�2~d�J�������xG�^7
���T��BlU@���yUX���Hм��@~&��9�d���cc�&�u/hº��#PQ���^�h��}ߨ�
�'���c�>:� rb�pv�Ns�ˍ�R ��<j>q?�gy��A��35���/�����S';3$�3n�
qН�,Ă���ƫ4���)Hxz��z�K���3p��-���[u0�+���EU��w�yuꔥ��y��YY��. �ן��t*�AH����&T� |{�tu4��b����"M��A��R��� ��N�D�T�hh �I��J�2o���>��Hg�c'�{����g�)����k<C�^5��v��ym^�5��h}$.5ժ���'�������i�/	j.�����ׯ���bHF�� �r�Q>�����
�t
i-��MV�(]X�n0�ls��`P/Nz�2�m�H�f;��Fl`�;x�z�3���U7�~�^'[E��\�#4lu�@�h˜s��`5 l�9�[�������ۨ =i&-Um;�����n�D.��W�954�T��r혝��(l�K�2�6 Se,���J�<| �b����t�Y���KG~w!8?o\�;��n.�,ڂ^o��e$��zk��i�Ĺ��, r���Blm�
j�ttH��vK���q� rE��N�{@��cӒa8��� ՌkFQ�� 0�q��:�	�����7s��N�Ϩ���b��S�d�Ǐ�ū[־�PS�C .�Ȼ{P�i|�8��DϿ�`�@�*���B����B'p��(ۏ@VzvJr���rXu0�#U�W5 tY�g��9�������U`ݻt���S}�����]��4+���Ȥp�:�_� ��L�����ޑ���B]�B

������I3��)Y�Yt�����]ɏ]��]�u�fr��,�w���|�O߈��<į�X�<���R�2��?x���pNE����z��
�P�4	]��>��mZ�Ȕ�}����L3A}��9��qS�D�`��O��g����
dĈ�p����b=KAi>�O��%��!le���xi�O;X��"s��s�����9[R8�SKՈ�FT�>�X8Fń�����2&&&<��˩��m����)6eA��	!�yD�ews�D����9�7��� �=a�'��Y�k�_��?�;̖���3j7SG��}S�G}?8�xX��WH��^��V�b1?|�m�q������'����Ĕ�B͊���{p���t��ԯTn��8*��I�}����(].Ǩ�A"~��Đ���ej��(=��"C3((n�<�����W�9S�M�e�����1���~�)��S�r��'�\}��\N���X��"=�Aq���9��_��n��J@`�@��CZZ��{6}E:q��
��G������u}��?��1��_�v0��P�j��t8��VSS������ 礯��v:T�欭@8��"�W�Ƈ��Y��s�7 �.LZ�MM�I�?~�G��1f,ժ��Oq����҉��D�Hr C0}�իW���s|j�+���,�eao�뾽ZV�
�q?�:���t7	 �� ڢ�� ��:�B�Q�u�~b�7kV�L���z7~N󱢧��VyVo�U��W�J����[���q2�u.�^"x*jZ����W���ª��r��k��>\�[�m������a��9�C��2`��9ن�&�g��2��֫U���q�_�-x4(�r-��_�gzx��蹏��Y6rKGē}�*���OV����u���MXQO���
��<|�]�8XY����?+����333K��I2������`֨<��WZ	L�ȴ�vi�]�����N�Q���Q$�~��;hsp�d/�[d��U�a��	{\��Yk�<���/bh�bw@O,�u�'�����~����m�ˣ�¶;���9Ѻ=�֐[���ζ/�]��+�/�p
k�g���Ө�D�a��v���h�3��D�9�^�� �<�MhN}|[[[7l�[V~��}�2z�s�n��Q쐘<1�m}��@AF�O�mV-��c6��u)`�Pk|��
>��߭J���A{g'�hj��N�[��s�<�.%̔UvS���EN������9=<"'}�B(�$ r֣�����)�i�(]m��A�J��m�����ʡH0˝�åa>B���>a�q>/�Ұ�J���B.�Kn�.M�f���d�+b���)��k|�O,��ciyyfQ��	�v�z_9 u�k��Ћ���D�n��K;�XlA��q}?K@�� KQ��G��|�+)Ͻ����!�Ƕ�D��c���j3o4���_�c/M���BT��]�gj��L��E�n}�2���~�ʂ������c��I*����a&ff�<;m�\\���PJ8.���^ ���б���@�-�Q�x�c���홚pb)~�K�z��\�VD���А�1a�=		���ʬ���Ǐ<*�~��
��y��s�6	�6K"��O�'&9�x \�F�MU�y\<��lW��SHL%���G�����P�!Q�k������@M�y�b��#'u�~���\'Ćv(�"�Ç��S��%E�g�k%#�L����Hvgr�	����O�87U��I#�9I��U�.�ەcX�5u����G��1�ѡn�L��S�F7���YI��c[��ј$���S���Zȣ��e>�,��SJ���ode���&k.�=qUܤL�*���@̖�%=�x���B[甽�օ�\���^��@:�L����0j֠�����e	*���hh9ҟh�s/4�J���z�4w�@�����'E����CD� '�#	������@տ�K�<~aՇ�+[uDL����ys--�ᑑ�I�Y���R�k��}t����h��L�ﺥє����S�(�s��4��Ż-HՒ96G&G��!���d�*d}�`e�`t�E���,��/��[z^:��=��J��}j�Y�yՂ<T���\�En[~(<�&B�V>-:Q�V��gb��m #��v�0��uZ%�h9�aXƘ�R�೻k%Y��e��^S���,��^���MO��سsi��T�4�����jA�9CEDHB)~�j�	�Π��F�ݣS��W�LL�@���9[�I�R<3��w�Ao���C7��ʹ������e%�<$+�F���J�hDC�A�(�)O:�G#�4�&���DscP�K4.R����x��hɄ��-��� �&(��@bdK�㭻'n+�n��gfbb^5��W��C<����Hs7�_�x�׳Cl�ǀMǑɊ��m������7�@�-/���'7�js$�������R�ݚ��l�6�k� ��f���S4�K2G���(��۩�],��UT��������:��_���h�#"��:���WF��� j.mr���!T,�R�Dp9�
;��*�u~�K#?��IQ�$��h���\KP��Qa��^s�V��a�����J����F��T��h<wqQZ�Qua���#��'��Z��WWW2��C�^�o3�-��=�����}m�@���.�Ǯ�����
�Ĳ�?�����x?zQ�M�CՀ��v5~�����&= mP^���~��/���Q�&&�A�X�1~����獚9ny��39j�9<Z�DMǸ8�E��׮hrݞ<W�u�	@I^��3j��y`m���xQ|Sm<G�#��&�ˆy����;��ƠW���,�wڨe��� ����H��o�&_�7py�y'����-Ѯ.1MeT/Y#����:�O�a)��	і�P5�\�&w@�H O�14LMi/�J�S�m��SļԽV&�brP4�&���Jnc륻Qa�E��_��-P�;�4��S5VxÍw����&�f�ϟ[�p� ����(kt���q<ּk�N��-PP��n/�����8-��}�ֿ7�u�86�0���~i��g�{��T�P�'�Ⓚ�A���9N�.%����U粹��UP�u6Q����k<�x�����C�
S�Qhܨ<��3)s�N�,F����gj@��� &(9�.��P�V;"ö��\�my��5A�
\��Y�ʙ�b4_)'�)N��(=�Ͳr&L}����SB��7���1��?�<�u�GM-�u���%���]. #%eCU=O���v�o��j��b kf�?�Vk�>I*�1{W�j��|���i���Z�a��<����B��%M���s��"��
?����vj,L6��
6Ѥ��Vrw3����Y]{hn`�Um<�;�Gu#�ɠu��Y��\8�F���ۏ�*���ɩ�S����|�Ԧ���N�FF�GƘ���kU�2lk/	�Qw_�"&�y��J%O���(����l���&��h��ut�(`'���h�v\-:"���i�/{�Uԯv��Q�`#�7rrrو�%n���X��K���|�]ȟH�p������s�h�����r��p�eP[���Z���&��	B7İ2�9����ke�* �p�Sm���)��yv���s��T8<۩Yz��eZ��� #���%#+;"@[�[�;%����LAT���6�SmJR<�kU	�b�ыss�v��Ҋ���e�5S�ˏ���S�p<����ohƾ"~�Tc�V9��k�b�O��	�5`pC������ӯ���0b����)�k�������᮵�S����q-����lg4�mNh7��
���9���^���LL������|���"�_K����� �"q �(��&�Y�;[юEA�ai{�V�)y��tvSc���`�Oh�(^�  ���nOU�"���G%�y�@.�ɣ&� ���@�̹������3mr�oy�� �l[�^��oAʻ��m�bgǻ����R��TU����Ͳ^�unp�XilCt��4�2��z�`n�2�90��a��/1)�0�
Iګl���iS�3u��l�7��$b2���J��LL[(Y�Y�o0�7֥� ��+Fvp S��#�EG����vK�{& ������WT��_eOOO+k�U���\���n�x��^+Y��On�]����� �x9�n LLLg�_��:����%Zsb&ʹ_��M�?<�;!�ڡ�����l���#�Ȍ: ���Vf��ǭ�e):P�F��S��P�c��5ǔ��i�(�h�R���tT�����ï�,uTU�+��^��� ��(\.�X�>�ӓC}���m ��U�EZ���c�N�Y܅]!A�9�B}dd����x���Y�`\)�������O���.=��({b�}8�%�2�_�@UM ���ר�%a���H��r��x�D)����a2�ȘQ�j��޲��ڳo ���[NԷ������UUU�t��ψKH���M����-������,m�e	Ү��������c,�`儺���-�Q���W2f���/��@�&/��ݞ�L� �%r�������\�������3�c|	���0��[ޣ�O�#�K�.dvﶊ�R8�86C�mh4l_�7J�l��%*]up}:�o��DR1�#�A��}�uƲr�p@��D��o�a4���Ȉo��^PSS�[�^P���Χ��{�N�&�5��M���s╁�$��kW�����P��9����U@ےS�Z�2y��]`���U���|(�����U��	�c",���^��������F{�P�,�ge��7�N����b�qxBa���O�ftۙ~
ٽm���g"���֞>}zv2e��A �
��г������9��wm��r�����vq��mC`l������D���N_H���������0$�~y�Pn�eY�]nt��AM����.%S銹5��m[��y�{i�K�p��c�E�xT����!��� (zg���~r������b�`6.Hr�	�ͷ�Ir�y��,����u�c�N�}��M���>g�o�U@����T���{�T4i���&�T����͹��b��9I^�� s�~B�٭�Y����>��3�vJq�y]g��ڟYtï��u�M�3���lN��m��uޞ'����<t��S�9*��K�	������mDc��X��a�@fҮ�;����!%�f��웥m�j!G��Ͱ\Qu��(�a�/��RVV֩�^x��������ބY��^*��sddd�I@��u�$�seY�B+��S���YV�a��L���l\%D**>�����xiʜ���l�Y;;���P�P쏋.�2<$+��}h2��t�$����U|���ð��pbR�h3��(�X���Owf�|Ny+U�����98���+z$\�Dϩ���l�0\��\u��=	^�h�W��9���͋x_�{��5Њ@�� J��ؑAUwOp��&�L���J!$tXkkk�)A�v�)�#
�"�;�+d����o�W�Jc�AK�]�����oy�׈IgbARp)�\vڟ�z�B+&�Zվ�ë�z��6���jT�3:e�{ssS���P��Aٰ�z���ÇWH?*�'���t��#d��o7j����P8���NVH�*YnRj/V;4,��!�J&	C��hb�s�v��1�g�*�P
'�&?� -.)�b�R��b���o12Y�[R���Y���|ө�3��yy���y��)%%|�7�J��d�L���&HoD����?A1Ǩ�!�`��eb\�{p����	Y(-m!������'�S�j����;9R:������}8�UO.�K�b�?���v��: *�l\��=1Ra��Y6���	tL����X咨�Hg!�DDB�	1]�%#6�̴&����MdY'L-ݯC%�����y����w���4��������Rn4�es��Hm����?d~���-e_'�Ǐ�H���6��lƵ���b��
W��~�u�޾҄� �XwjZ�����'ۤ��Fz�YO����a)�7�惰�L�:1z��u��"M�G!� YP�� '�Y��hV�B/Qx~�W-���BFA1� N�9��l3`�?ˡ�;W�z��I�N�p2[(�R,�G��}o��U�]xt�-s���X�x�.��J߈��ٯƤ��0�E
YW	�19��mk�j�em��as�1�����x�~~~��m���#.�5��ԯ��S7�Jp��v�sxdhC2��c��sJ5�{����.�X-z�I�P>��лߖ�"���b�BT�b�Y��F	N�VH �L�|ѿx!���dB�ExD����lc6�2�̾ք�E�HrAb����qi}i�!��(�����2�Y��/��YH��I�umi5�o�_N�(J�XTTTɥ��#��s��Tzg!e�n-�(�Y�����TPP�/���,�C��i��-��Ŭ��;,�fxH���mS=��D���2`#J����is�8D}n:#�7a-������@�6?�W���U?�O�X\'#)99�X���_5\�u���D�����++�g$���1�p_��;n�h#j!)k3jsڪ,�|�g�@,}���Y����D����f����"�9����y�# �r���hh �{{ۀ>q���XP�:��T����zaw[XX�k������N|�>+�M��~B-$,Lq��=��n�8���/���b�`�`	�m_~ä�x�ڗ�N��
��""����,Uu��$�^�f�]=��߯R��y<�]�E@=�Ĝ�<����-`Yb��8j~���ܱT�pV>����/`�:�2��=��ػ�_�E<	u6b#�C��O������?,D���	(���*7�0z����鵡v�-�>+@?G��~���N�������������o���*�V���Q �:z���̌�w��D�����#��J+u�i��cbff�q���lc���=44�~�u8-�iJ��/�O�d�^]�3&&��k)
���@%pmܝ����?9*��0�fd%v}n������>A�EX�m 2�hlP�BOQZ�W��>*���N�����G��)�
��A��cbX˥��ED�2|/,���6��\��Mr��� /���"�e�L�.�R�� >S��B��RgT�I��!�CA�MǪ������y�� ������t9Zނ"����}}��\xnϱ�pp����O?ݞ
)��O�1_���?^ώ5F�ܞ�NÞ���Ha�N~%��9� � \��,i4Ó�K������M�J���N$	wI��GX4}��[e�aC]�#G%%������۪�L�Rrb�y3bc��r�r���V��[G���,T=v@Ѯ�Tť/�z��V��#�����fเ��a]�Qk�ql\܂F�os�h�Ġ�����*u��6,��%F� ��b����4^�2����E�r��q�����'ۅ3��1�7k鴹�I?䬤�ְ�����D���{l����'���r$�\�-�A��GU��3���4L����� /��_��;::�X%!~��p�������g)��7�qg����s��LDE�X}K����1��1/$pg'�;��HD�ۼ����H�ix�|q��O@)��px{WW���	��o9_ǌc 9�1(Ր�
7���d��j��HyQ�7�<=��q�9[(W��{�����Bt�#D������Į!0�1 dL�M��YrZZ�>'����?p��'�g��i�'?'���G1(�<��#���\�������$<gn�1�N������'V@mw ׽�=^%���;E������),	�e��j�k�b��~:���� T��@@`�/`�ģ�9��xu�AC⇛�$''�%#�S�9ӆ
"Q���������ڑ��2�CF�L��iv�h�5a��҆��@�mw�((v?y	����g\�����ҩ��wc�UHӸ0/�5^1��W���g����V�B؏�ѧQ����hخ�M(h��ֆHy��U��z>��GGBB�{T���t�g80KQQ�0�jX�Ǡ�`���4�cE�+.4�[K3ns�ק���m�>~�_��2�6O����۳����c����x�p���'����U�XB	��6n�Gb�J�#gm<�UVV&-�))Yu���=�!YW������Ԣ�S�f1����zW�͛������5Z d������y�D�~�F�b5���Ѐ��(݉m�d������;���U��8뾄e����>�hC|ZZC@�:����`2�B{-(P�R/M��4��D�qJ���,,r"<:��O_F-; 8�.;i8T��DEY�&G6˖���[`���5*����P}�*yѽ���OK�o���pu�E����wDԅ�hZ�,9999,�" n�����_���6��'+�&V��� 

N�z�28�		���j���K��5�����0=�}�����͜�$�ಞ�j@�f� �Hɜ^.�0���|r �4�芒֢����zyy�!��Ć�� U�U�f1L-p������F�=%?�8��v�;HQ7�ӷr�������*K߭�p��4� f��p"��	^��{�-7f�y�@J]�ޡ���V$����iEh�x�������������D���$"2�=��r$�p����4��H�S�2,�����'-�ИQUU�l�}��ʫ�9Y����ER�~:Z�
u�U w�'�]DD��b���"��0`��0�5���3>ˊ���	�n���P; X��f�벉��s�X��N(���sn���d&���[�Z�y��ĄT��� �F��Dܜ�q�������7��J��Ծ\V�ܴ��0O?��'H�(o�����bwX�Z���a�*m�h҂�o�b���ZܶM󳋜�V=>IK#թu����;J��m5�$����Tm��h�
�H��[����E��kn��N�ONN�.2۽��<iѨ��:���ҟp	�Vơ�8@W�4��l"�0�� ��%���+GJ4M�;�P��]�K���1z���� p�r��{zz��Irߦ�%���z�����:��M�c_&b�Z��HجƘl�K�id	R�;ε��T�aP�}k�Z�ι�HU�9�`���a�-�[, [
�=$�˭��
M�gb��a���+�rQp_� �7���z?C/��9��]�P0�i����<�-,<���]ㇽ���Swo�E/K�c�	��?<�jzZ��>9�h$l������9>@��wF�E��"�?��^Q��ub]�]]�IE�h�Aokk+��/N�z�Ѯ5�U�^%0���z�)>��[�bۗi�1����G������t��a�Zն��o)`MkZ[['�;&����>7A]�qTR��;�;~���< w�6���������Q��M/ r���|��hDQ�f�6&����]���k/���{+��Fܔ�x���R�Ԗ��G@�BT�\�u
0zP�����Iݍߊ�>:*h�i��Nfbb��}�y^.��L�������穓��%P�P�?v��`T�,F i�?sZ���}�_ѳ��G-�����BS�uS��ךR�x꟟-�T��e+�i�s�LL��0ʖ��y��A�a�}`А�b�t�3���(�O_���Qc##bi/tJ�Ĥ6�^��2C1�����^'w}����g������%��x�Ǥ�� ��A���=�}
f����˗/�b�3��cf����?}5�%�^�fؗ���9G�&�obc8��o߾��Y�����@YcZ�7/K�t��!�:img��k�~FFϡ�����M .�6
�iEFFf3�Ɖ$��ȵ܌�~P�Yq?�ێe�������|�U�V|�����t�5}���ۮ���j2��`nY�\H$�k�̠XB/{����W���3��ଯ�'\���RwI���s�&�^�ޜ�>�	���́'d� �6z�bVt���V�ii?��А��na��#mUj0u}��_�~�<�Si�!�����`�5���뎶��\_�B�����8���[N������/k�2�����ϊ��r�M5���ӿ�RI|K�ȍo~@���f�A��F�KBB�ԭ�d��_ݘ�W�p]�Ԭf�R0(��O(ũ���ޱx�>��#�^�ux$��4�b�h���b����J�ۗ	2�!�iל� E���Q�����0<�lt��2�Z��E��ю0RQ�xer{-�dڠ@V�{�"yN��.�+�qqJ㖕c*�J!�N�PB���s�Xv�9Qh�n���� >�>����hUb�~fZ����Q�$,4��o��X}u)F**�:O��ʍ��4y���1 ܳW94�?�q�qZ��j�������KBf� �3rD�}��@0�kV�~0�I�DM��<j)��F8<<���?���.���1� x����*Rͷ7����O@%� �Q9���P�룢����M8��#�s�)y� � �!$���XM�Y�6�51���e��2�0`qII�_�R'��BO49ͰH��UU�A4qHH"�w���edd~Bhy8p�����4p�;��R_q[�t�૙���!��Ͻ�E���������KU/.�����!!�.*{�F�&N�=����"r;��WU]#3#�Y+�]�7�}����=�KJTz}���t�OO��}fO}2(2E�'qQ�$ss�b=
	�/�",���:����}�'�KE
_Bࠛ�[J( $���Qy����=��J�q��N,���*�ά��xy�.w��|S��R�1#dr��u�]IH�m������Bq�]u�]��V��Y=���"$$,��
��²��}��,]!GKpr<�>ܞ/}��=�����ֿ����CW�>/ח��ϣ	�!������\�ܐx�b��f[�(
v��زF,,8��WC;��W�5*u���'跢	�!5,3��9I�(M׹<��������↟<����$J�']!��������[^D'x3k&/�n�����i%�t^S +����]��G*Œ(F�I�Vg���π���e�iE:�5^��^��7����8�˨�ѭ�m�#��3��R�
3�7�ޠv,��l<q�tk����!%�ّ�y��%���[���0g���S/jd>6��y��݃7�`L/Yt�]��-��wŭ|8��a	���9;�n�F���,)=��L��iq��ui�ŋ�����?����x6�������_�QK��onN�cX}�#��%�h�t��m���m�K��T�Eaa��FA�^��/����V�A������ӗ@S�����d���*ɔy�5T�"��d�2��.B�kLH!dJ�d�<�y�K��������׻Z���s�~��|���9�#<�R&�=�/�42�]Q#m��ֆk����z0��Bn�y� �V1�d��÷�f��g#��'\��������)R��q�ƍ�;�7�:}1KNXLT�yS��3d-��o7���[��Rܰ6É�����:���1J؏�V��l������R��<��F�v��LSGdRh���)�����=�X�P����S���c���C�{�2�����hCb�r�ߊ�A��=�Ol�OA�V�[J��#l��Q  qߴzJ��#k����	�v��LKS�g�N�ph5�~������K�����c���R%��m����-�3�cʿ�K�cà���sM�]M�_͚u��:������h���ջR	f�w��&~~쑑�/�ӑw�(�C�/|� &a�jZqk�qj\p��h6�"�GR�GN��p#O��m����:�.���+說�֢"�uB�'O(�6b6�8��_2����$�y=��V���{�|�Y��j��������9��ӂI7)�x�ˍ���g�_L���3���V[[�W�f�>���&!�9�K?G�qsS$1)�\0$on�I
��U��6�4��3�Ju�u9��������>t0|+g|�:��U!�����p�J��5�5�n+��t��/1��K!K*��y��z�PY�_0h�	7���
��=�.�����K��]<PRV\Xxy��<j������tp�Nݎܧ�ϧ}_�^�����>Ur�Y�+ �����f���v>'{7]x�����iZ�3�d!q�P�w]QY�Ɗ|Yľ+6�z�C�������c��݊�2�����w����Π�Ҵr�r�[�C�B-^9y�5��Z�������F�22u���1Q��}+���A0:����ECְ�S02QЗ�tU�����-8S* 0jc@NK��S��t��r��8[R^޼��F_�'\�,��d�R-l�Be	���/n���d�^G��a�ժ��_J�fج<W)4�5s�~�:�3L�b���7���~n���g��)E��[��ȈF�$�9U��xbp�г�Ҵ8�!���&a+4څ(��!�����Y^��󴴮g�2��d��
׽j��5����h�o����Ce�܃�ß;:��/>�\�.�Hi�4,�fE��	H�	���б-�АX��� ͣ�ZOGVB�f�;pB��� Hf�&T$��H�M�[��t�򜂬��La
��]��L��A։$��O<~,<��t�-��-�ZCY���l�<�춴48K���*���KgfZZ|�,V�Ab,&���ꔊ��H�|rہ����������WJ�K���d�s<d�������ٽС+dAIm'�^7r�C�y��>@�վ�Lx///O���������W(�JO�5ae��^��7���L.A�>���v����ZH�`1�;����P�f�h�"��S��i�%�6(my"�Z��b���t���i��R�� ��	q��"���}���m5=���ޫsy޲�_����D���?�,��s�Q�*�p��5rޣƊ��Y�T7)ף|��zn�^�54�E(�#����l���C#�͕9i�-$�PY��=H�	a�˯��Q�v�&%a|�SEN���w�� ȩ�X[��\#�����A�A9:p������[�Md`�P������)����yP&��8��M��L��x~M��\v��~��+�*
[}|#��Z/Y��U	��&���C1f�w�"9�Kᔃ���~f�F�UZZ�\l�H�,�%�w��$q�"�꾉�� ű��d\b��ow��%���,y����킾��XRbi��8�S�1'�*.iü���v����ZP�R2�3�ɈL�v�MK9�P���cv "�X�al��Ȑ����h�H���>�`�����Œ�{�.C碕-^
�0c`ijg_�3��;	�����Ni7vu=�����ӄX� p�^����˵���UG��炻���ѐ���ʑ�a��T@�A��y�e��(�-
K��ө1�w�6/�)O%##s����,~d�|���>��Y�A�Ӏ~\p�lWi�"��E�%'_j�#��;��,*zZ�����<P*���A-jA�3��`R�Ix*i��W����<﫪�aV{����0���ןC���)�.�J��꾀52H�`ς0g�����Kѿ��}}w����A���P�*�")&�l��@ax��)}թ��߸c&��w����k���|Ԯ\�$B�
 ��� ��]� �(���ɉ��������ƵLv�IBP�6U��%:Rv)Z��:R�����'K�lA?��,��m~�Aua»-���͋�m�E����A��̘�.�"9*���Vة ������H^U_��u��GJ����,*�[����\��8�\\ L��A���l�dD�����/l}���\�[���an����||XaX�.]�cF�47 ~��@�?�ԁ<W�y������D�ټ�
)Z�s0a����T��Řb  � ����ս�}`w��.,�lGT��_&'wW?C��Eí��ш&�����	z p�J�m~K����?&qk>|㛉���5Gv-�����H���H���`�^w�/�&i��y����Nj�k�s����1����D�+$�zuۀ0��<�A"���G�k
?�P�9ȹ���C�)���yDb��_�u� �͓�0���;�>o��x�N3
*�t�C���G��g���~�����V��h�����N��CK#��y�bF��{K"ș*S!&�U~<n���ݶ�+����[.�F��cb�}�j�5.�ݶG_��e���"vY�;��9"+��Τ�f�i(��%<$�ur�Ɛ/�������HE+��F�����b�g�gz�G��n������������_Q��@j0����>_^E_��`���zT:��2�HIJ���q��ܭ���?�s�'�L�I4B��cu�6$} OQY��41f:��e�&9�$�����4��'��1�����{����D��R�>�J�k��G�
G�=�!`�*A����1����`����u�B>k5BW�����~�W���� ��<�����+	7�ԅ��;�k�=F�)K
���G�����(D�n6�-��޻�HUݨT���% ����B"ӭ2�[���~5pEe�&%L0�Z���j����+�#���4=�|%�� z:ܚw�żX/�uD��X!Q�B�*�w
�
�m~��Ǖ#��e3&�h"d�zvn.��ӕ��?�Ԩ��
��5�Β��<Fጞ.樗/_N�"X�|�n��s�����p�r�Υ�����zЇ�
;?����5�}l������Gѵ`B㚦~��kt�ʹ�8��ӌF�z2{���~�n�����h�iK�<8@���混��|h���U��M�B;��4����0ԎeС�E����ڝ��-(߿�%*!H���ku����h�ǌ��̠9�����#���)��
�E�N�;s�UJ��9�Ԧ�����[�=�BL�[�ѵ����0�`�n� ��Y����$?�ȸ�'Lο�x��P��>D�]���	���=ZbiJ1-Z
RZ����v��Uf����W������%Y/+��l�����B.�!��?6�����)p����o��$�WI�Y#��;W��o��X�u�Lo`^T��b-ww�$Na�@{SB�=kmmM4�?�`�����$!5x�=��Z[^vy+p����+b�kvnzz�ka�9�6o��}Av{�D�����n�n�k� �b����n��L�-!1!%EN��D7T�8j��/4P�Yz�״���'lɃ �-)&��kO������1��(1��A����X�"#bPr>\������ߗŖ�9����W����&M�L��bL�-���F���öN������Z0Ů&6������9ڠ(T���?
u�(��{�\��*�㹷��l.Ҹ���������k��K�L�o��G��ۑ��е��ފ�U��x*( DbJ{hNNN���H�F��Ɲs+n�-6�;��kյ�v�gϞ9ܔ��OjCZE�-��ۆ�:���(H���f�i�RǷ�7�0�E�8�"����A�@k�����F��ZuSl���.*��N��n�����ǼU&��K���O�C����U��q5O����ȹJ}��x�7��~��*�'���S�>�#Jy<V�T\��g,��weIU�zYXNZ�
	1Qx۹�8�T=�5鶹��a�j�,-�1�1 x\xߘJk�����E)�p��3N-�"�R �'�A�qf�\L��mn˚�
�5�� ƀ5x�A�#�����#/�Ǎ�X��gw����BTw��Ϸ��i<|O�_��o�pa�<��<J����>����/�Y�qe!�Ƴ]�q�H���s~�$��ƕԖy_ `o�a~߂�PJ�������h����-��C�X�6մ�jۗ�/ԅ��fټ�M�|�VD��v11)i#��O�IC��������p�y�}��O�Fc��~�A?�@�����h���M,,Nٞ�?�x�모h=m6hC�<���.J2�~=��E�4U��W���B��#	�dl��t�������_��ʫŰ�_YwFS~�T�p����xʎ���(6O?�e�;0N�JR<Q�	m0����ur{ �>[��}<j*R�dE�x����-P�bok.��pr��y�g�M䝣=%��|�ʴ��ߚ�S*V>���.�����`����*�۳VKKW�	E�h�@�"�;Kк���� ��W$JC�����cv�����n3��tէ��	�[ec��N��^��oŷ����ݛ"����ի�k��+O@�c�(>/����&�}�*���i)y�Bw:�v}`v�����K�D���Ŷ�葦������B�l��b���W~����m�$�ѝ����'g��)8:?��n�i�m�#ˮ��{�	��ĤKf�O��t΍�����P���,>��q�6ԯ��e��s��_�u[��g�ׂ��Tji�P��#�	>�}�:׿�&#p�4���n���<���	����1�}��O�>�����<����83��9��{��o��,:���V�s��cY�@�ٝ^E�R��z�7�O��o�]�Md-�-{-$�P�4?����9t�2Z'w}�!��\���	}�}����ܗ]��`�Z,Ō�7x����u��U焆{S�;���`*�d��޽�&���#��|6��0`���P��kH�A =���U6�e�a��ﾛ���
��g�N����Y�h6n���fC���G�be��D�m��+�f�%�}+�qyIF*ME��{�`u���u.Ļ�Ľ��y@A����*��W��-zBJ�B��9SnѲi��ɲ�S.��%Lx�����t�º���2�];:�ϐ0Z;���K`V��pc�J��Uˎ|[pe�r�[�<ܝ�h�&�n�W��-��Y3RN#�᫪U���iŘ�V6I�e;P��bifO���~�s]�}��%�s�\0,�B8#~:k����"+��R�/md3ML�?��!Ѳ[M���p����<��e�9\��'ʰK2;�g}&G���_�!Z�Ko/C��@��#���*8�k\��^/ ��`�U'����,�� Brʩjҭ�31u����ܱd@�^�_����^���b̔W�1�����
���r��D�1�)�_�:���w���u���X�l�|Od�"�����i/\B3#����м�^\���f�E6A���{W)�xM���#����O����}g�D1��g	���1�t��+�Ɖ�� 	��'��x��L���6MM� �b�	L3�T������[�b�XB{Ԟ�5,n���gx�t0���ߣ��v��P31faqqR\�#/�T�r�n���Jj��~�;�>�͒3S󨗩��8�F&�%�m�B�k�@	 �S,��ڊ� �20�KkJ�/��:��LCI�g�9�Y��k��쑽SWU~_�͒n pF1����z�{iɮ��T����[���Iե�g��[�#{�2�T n���J�!��bV�=�ťw��TUU�$--A���no����|56�+�����2o��RO~�q��!�	[����AʴЈn�/�[s�K�����M|�8h��V��w��E�"�
V��Tj�5����Y^q		-��C!�I���%�\s���*߰��=Z��PÌS����I7��P[��<����0.{0��+^�MZcj(%�4�bXS���;�s�ܷz�(�pи[UEq<�+nMK��.n%�P�*0��±��?��81��xS3~��ɝ��xZ�R�RN.�R,b �c�{�-_AL��k��ڟC?�.�g"�8����3nx4\^�
#�(�)s��cn����yb�s	���&���#��W߽�����:H>C2Ԩ�


%g�c10����\۽�	���C����;��^|���e�X�1/>s!T<p:�%�0�kXkX\P�X�wk�{�tA��h�.��"���'����̐S/�;���,�M�J44d$�m���\�e�C}!k\b�Od�?U鱓�L:U�b��h�l}Ae��;^��GV�!rSS�����E�M@u�m��WإG\�7��P�Rs ��������g��u����7FԢ����9���+�w�ueF�]�� ����t�ҥ?�����.=\nQ$'�I�N����b/�^҂�j4���L�hϻ�V��F_��ᑜ��{�[�HӲ�6�u���G�G��N��BD��?��L�&)|�Wm�:O�̌�i�P� ���Dpj۶Wϣ��v�����)�Y3��ΫPWY<EE0iz�}ѦՔ
o�CX�d#��Y[��[ь���_Wm]>�]=;�	~!����<K����:���kP����*}id�7��#��%&
"eiJR�j���N�p]]]�y걯��! �C���^z�kx�`�T\��2o+B����gMӓf�&!�e��Ԟ"QR]���f"*؍T{�bn��p��l�`��7%��M8�筦T��\PL�g�\�QY���c�e\4d�2��%��J����y�n����w�����ֵ��a��G�'���R8�@`��Y�U3dq�,!�C?ґ�\YBk=m�V�g.[D�{���X�C��O�9/��a�9�ɍ���_#!"$
@6�.�ٚ0-�㥩s�yWt.�yWTd��oؚ�Ԝ��b��򑢥|m\���kkg�ք,'Ǆ/FtJ�S��D�5ł��k����x	fmu�*����x���$X��(P�^'Kz�P����,��'�+D�i��Y����*�p�3y��~P�0�@���q��Ρ΋f�Fu%%��go���:R�C1��w�u[����l�p�Y+W���h�6e`�ڗ�Yݖ�q{��ʩ��')�˗��,5ى1C�2����j1|�v�;�
�)�� �h`�LE��c(h�Z�v��ګk�]��~ةT�!Ǡ�o��|�9�rhi˻��n� �F��E���{��Ab[Ma~��&��*r�f7J-�VB��qݫ����,##-b�;l�M\\^�B��磔j�ni�Q�=�)p�n?�(�
��l8�w���x8���)��T�ST�Q&
ďDH�vx�ܶ/�מ�=B�sA�3�N'���Ҽ�|�b��H���1� ;� �3�'�&���yIO�ڰ�1�6�u}�p�b��&���$�jv�⿭}n`q_�@�TLn�M& ���)K��bd���Jy��!�d��Kx(��s���ysNR�"�:���O!G��s�0ސ4�b�9�_�ܑt����������E
nh�e)F���;��@�=�T>d��phHj�����y'��xJRm���?uj[ ���Γ��J4�[�B���Ş����:��PȽ/��$���r
`������)���b�9�^��~A�fsh�"q�I��cԖD,կZ$vtvf�`�(�Y�����ٛIo�QYn i@Y!�*d߶�`
3��d
��TՄ��e$�ǿ|�N����d�e�~�P��m\	�<�w��.�9��:4��Ǐ��'��y�����D.�8�X�b-�y�|�&����p�ʯϓ��(�!� zb�����,Z�vX���<T�qg�[�A 6�ef�S@@��2���4hrP�~���$<��@O���'߸��[�����ZE��4�Ȍ�9�<�h�l�}��mi������|zq�:���9�F?:���\N�}��݅Nc&2�.%��)S�����{1d��̟_{ �0*�4�׽���� (����~O���n�a�y����C�ޔ�f��'&��������]٣�ο�cc�sB8J.��Ӏ,�LE�-�}�:;;�<��0d���s�^~`�˃b��
�eJ��|���G�#���׃ɭ���X��G��>B�eW�3P���L�w���k�(��K�w.n4j �Z5�>��-���F�i�3)(����$Jظo�À\����VGG�L�OX��F�bՏw-�4~惠��~�L[����SBH@U��Cw��N!��Pz�������.�sD�͟?խ�\�[�t(q0q����+-i[6 ��>y��h/4,�R������Z��-��+F�% ���*%��݅|���O�UN'4e7H����2 ����$#����j�?���R��\t�ߴ��/�B-���>@�P3(5VYn��Qk���Z����;�B{߂�^�,;cE"���9��^d�����pt{k�YQ��Bs'k��[9��?ڈ� �/+��p�|�4�/�u[l����s48޺�� 5�nB�*"Y#��nX8{٬cA>ˡ�<�-��
���|+�%ed��\T;���L)TiF�˗`L���\���N�|���W�L���B�躴�����7U��3����!Yȵ���V$"��$���(e����(�����E&���F�ȼ���J�Jޚ|��dO"}K����Xihh|4+��s���Ы���������9U�i�����������pJ�9�'�� '`x����#�ED���m��Մ�$�_Y�5�YX��v�	فʠf�aº��}�p����9�R����^mv��imx�&k���}n�91�>����6/[��2��ӧw��x j���U�YfH�Z�Yn]:`٣[��8��t�,*j%�dʨ�h�{=���n2�J`�CB	��NAD����
�˯�����#m�ޘ��,ʊS����n.,/���Ȝ�y�"���F��t��`���i�2���$�� ���U�_�X$���1q<��6-��A��{=---;l+6Eo
��P��t�o�s�i�d�$gӥ�%�yߧ����T���B�p4rRU�����Y'�-����6�ͫ�zzzP������r�_�z�%��]�G�&j����s��3���pcp`�(P��D�XE����1S�d';���<t��4*ZKN��;µ����.�%�)��җ_���.��t*:>��![T��R��T�H�su��`�򞓪dw7 x~ʃ�������B��Q";8E��^F���G^�pf�ٕ4]�������(�#J���к�T�]��8+��9q�k_G�5�۲��b�d��F�9p ��\CS�ɸ�����H4
H����yȼ,�`!l��ۚ/�F�q��<�+�=�6W��Ľl��J�%B%�R�}���]§R��=������#G�qT~��f�RY�Ã��ș
fN��j�0̓��`�ُ�v�AN5�~MM�h���[�mi����:j5����H��u�1e�I�3�;���t2\����bɐ?�c*�9�
Nwg̝�eٰ�����s�|D˦��ּ��-���6�	��_O	�H�g�,�>���"��b��2��vB�a~����\rFG�������mn�KŴ4�<t���T�O �L`K7p�X��bZ���������u�
1�a������b?d�WTT<o���:UkX��\�G��!�W�F)��f��R"d�	�Q���([P:��s��a�A��?�c�}�ռ�x���`H ������K�ʲ!:-L]ީ=O��j%_P�y��k�8�ªrpXl(���C��u�Z���ML���xTv�׀�& ��ƌ~��� _=�Bߗ�:M��`EV�X�P(f����׷e��b5��g���^�,7x>C��nGt����7S���s�����;|�˘YX��ȃ���!�D�:��[�� �@��K�x� Ct�-���$Ci�Kg*?Ѓ1�W������&Rx/��ϣRڍ���,��u
ns�w��|pɳ.�X(�Ug���G ���v�I��65#����F8==M�|h� � �e|1?hap�M�W�4�WL��
��6��v���H22�6X�<S\+�ٳgA>�G�iե��_�+#���� �ʯ��T���Q0�T��K WWkwW�r�Pէ��uO�J@�+r��|?^�	9��1`�����7��BtCg}գz�î�d�WM9����-����/s0��M���l �Ƀ��qo4'M�?tВ�Ǡѯq '��s?����H���!�f����ɥ�
S^��s��8	�]�U�5>j)��	���U�M{��� �L׊ܫD����
u��S�3�t��X�g��F�����v�iOg��.H5	��k�]����Ǉ�Fa��`�UUR0`��E\i2���  u��!`8��w�츩�#U��O�y�_s��w؛M�2A)8�}���:᝝����8m���J���:@�����'űf�-y�hT������Aw��V�ŕ;@�+���3)�֤?�gP�Dş� j�%)]13c�˔����0���L�C����v���@�./4A���\�tG��l��N&��T�,
S���Q�0�ɞ�C�)�/��{8�@�,�ݏ�C�o�!l�;�!�����N[��O^K�չ(���pO�Xk5�	���N�p��I��)�N��#�c@I����ȴl(1&2��~�3��MT�"rH�b�:cZ��
���ب�G��^�~��`\ 
����L@>���V@P�B�:����>M�<(��;�L]5��=\�V���!!!ܮ�Ԥ�MǨ� I�h����Yaaa����*,��Zp3k������e��E�*�!G��ឫ���l8N2�#��;L�����g����U� )z�� w[�,����(&������a��z͑W�+++�ň��L��􇹔?�
	W�0	�)Q�b��Tqq���:0|�/k��?LE綐���K��ZlX��1����Ga���?�H<!�b��'N��V|��K3�?��h5@��hw��-�?ձC��Fs'�=~���Ϻ|�aN�@[��̏T@�s����� p<ܡ�9�����P�b������Ky������\�s3�'�}ǸlYR5{�P�H��i�*�9�{��$o��)ԪLh3�q�+|>I]­�$k<<m� ��4�v�ٮے�^����w@>������ ���ڈ�}��-G5��n���t��k��G(V\B�&�w	M����i����%(��nnnz�ǩ����th9�2��=�1�������C� �r%��,;�t��qWk1f�ݢ�.#6�i�ݼ�?|���pU�i����J�o�/_� Ou-�#�?8�n��A����X�j�YO\\��j���`�l���"q<J4$psR���:Z�)�U�뵡ؽ�,��zz��2�x+�t:�����)��������N3u��6���qF���� J�s;���?�Օ�.*�s��Y0b��Y�X�9(;W�BXcX��W�M� S� ?���{km_+�L,��o���·��z;,6�Kxo�+�ʽ_qh1|[Mc�}M]|-3�C��x�����w�:�,��ٸ�nLZ�>F�3 9���BY���0E�2Q�B��{���~[�{�h3Cڍ���t.��\\$�ce]�b	��mP�O��ﭞI��J�}dgo��ҡE���Y��S���-vX���_GZK)�h���V��G�񮒸G@���-��A�r�>}�*���H����sk�-<+/�Vv�ǹ� �$-~��Czi����e�����[�c�n��_M�j�?K�Ji�XC���&'x�\����d����~r��ꐡ��73�|	��	�w�V��W��-����!M���t?%�2����vs�}�D9�r}A��Nn*&K�b�}*�2�,U���6�
�r��֡sD˴w����VӠf�@hC���YTz`,k�L;H�Ǘ��w�z���P�¥w��<�>�+3�ީ��R	��vvȩ�0���S{�BMpf����������8��n5�������J����p%������9?�ك�/���Y�z�{��Gj�݊BL��ee2�{�W�%������黖��>� �z_Q�6�
ޗ��e�
:x&*��Td�����>>��I=�����}�ɹ��]��ι�� W��m����V�-eUU��h�1d���Y��NN������2ҡK��i^���hKR�5Q̡ՠ���^ZFN!����S�z�9�n���f9��d�ni?�Q4��W�KS�c>������Hb�\�&���D��۲�;PB��s��N�����di5����Եw|������^?Yi4z>2>���Կ�.\��o�#���	8U�J_I���� �
�����{g��@�G��5B�T��%���
��f2�m�ۓ&Q���鱫��f��y���7R
��8LK��|�C��~v2��B�%���!# :I#��;�I����Ԥ�G�ɂ���v�Fc;��t0��}?p���a3�n`�.��F����kj���Ύ�wr{`��8i&+>q9���n���?LuƐ4�4�IVR��Y�Wy��Xh��KH6�߷���fg�Fi�t\��Oo����DN�Ȱ��|��� ���Z+�$ɺ8q����D�௼$SWL��]t(Rp��� +��z@%��\>�8)�ռ�r��C?�⿖hVn�S��*��"����[i-�L�ּ�x񷗜�ж� �6}�����D0�у�G���Y�=C$��8�*
ep�\���e�gh�����5Ըu�DY��L�����)��2S�p���_�z�-�BX�ۙ/ᮻ,�x�PY��l�~z�&�KzW�u�~QbL[��͌)��ז��^�p/�=a����ϡ@t���iXt��I�Ze�<>�b+>RW�?��B�Ŗ�[dT�>������k��P�"�h�d�ʮ}A@{_�],ip��a�񛴗���ؾ�8E0�ٸY�����!k����3�c�òY�����FFF>:N��b�?.�ڣ(��xì��|.Ls8�fz�4��-݀���	Kʥ�!۳�E�7���������������H�5�ʇl���Ż��#�b�R���iH�_���b.r��br�Qp=���8�A�[����8�BS��b��c�d�U�Aֵ
�p���'��?Ys`�"=��(,'7V��2����s�����M��e��k|~$��I
�ahi�כWj]��3�l���AQ�ۣ�s�rf�����e�=�d��nax�,�zsGGG��X{�:@/��[�Tr�8۰x��G��km���Ek%�)f����mƧO���I�����_�#�� U�$��/@Vv,�a:�S���]�v���/&�����柘�ҤUђ+3,@V��y�q5OV��]��R�lȶ�y�w̦���n"��
XU�%V:�w�0d���=��Pk.2LZ��G��a�E�Ӻ>7^�֐�r��x`ds�����2z!���q�x/��Zzq��uu5���FK*�;��6	7N��9��/��7]����k�|t���_�G����c'H�WXxY:�� �9ӕ�t=NHT�,_�w����=>u�ve!t�$���L�$k0��5�F�s�W�BT�
�	�dIy���&��	@;�Voҍ�8/��>��ُ��<��֔'���F&��0���Ofw���,h�{Yn1(� ѫ�i�{=p.��*=�{�ɥ�R8�{>�"f�%��b,�C�{	��y�Ω�]ܞ��ϟt &��-A]bU�S?
OZ�3��84?:���ΨW2H`�p��R��mE}�=���ؽ���n��� �kk�<d;��=T�i����.��c��/[���W��`|��[��<����>^:��öL�a�e���.W �S��>��\ԟ�:����A��ׯ_'�v�o�v�^�#Ij;Q?1���!o|��6���
���GX��b\���0�����ŀW�j��o2�fq�c��+ip��K#����S�!p�#�6���G{q�f]�dI���I ����cs�
H����?��q@dz��9<J��_�K�0�b�`I������B'@� �]�q�?�{��|!�e�iIQ��|���Egk��[�7"�|��K⢌����Y�1�ʺ:���NU�?�u�.; "�	L��z�Ox<g�E]!!"��o��(��TTV҆�'�jh�R�z� %�5�K����q�ffm_{��������s�U���3]>`(�[��/ba��m3'ͬl�J���Wf֖�"岄�<��d]�
���gh@�ܬTM3NV���TWF*�,�gI�~�R��6HN�yP��F��s[�C��(��z�5cF>��w�v���k*�'-�3NR����>RݧȂ$r���[on��U���/�}��YÌ�Ƭ ��jv��������e>O����������2>���;of*�S�u������X[��p�����\�[��K�pO� �V��3�$ ��܏p�u�$p�������ȓ��r'��[s����S�:1�w�u��]���'ud�f���8��މ#o�m�V7�?�I�3..G�v���9}f��}���gׄ�s��jb���BC�Y<-w(����翍���˖�2�ӱ�ı3z���+��#��UU� Rfo���z��]�
�|�<���~8�֥�z�t�H�^N����MX��m��"���2�R�1a�}�V;����7Z��"]��P)))�55,�cZMM���U��N�>~f\�/a7:uP�r���ypo����jm(���^^ެ4��_+��QQ�3m�\e�I������:�8}9<�}��A�%��"|x��h�`a�fNN����i��L[������75Ȼ������S�Lb8��;ZZZNu<~:5�8���y�����77E�9sW�c�jxhGnZ����ж�.t�m��|�tȶez`s�C�J�����hm]]ݬ4r��]_SSt\k��z�Dqqq�Ǐ��쌌��??����7��~k�U���#y#e�R_���/	7r�?��:;;�VT�޹sGDL�aS#�?��@/��9t�E�Ћ燆���
��u"�5s{�%#�R���Iź-�?��V�ă�J�ȳ!L&&�����ٱccc�-H'e�}�toe�~~�^ѷ�EuQ��K��q2��ے����Ui����HH0�Ş=���<9}��g�9�_��`�?��H�j�Ib��h����P��y`a���p³�##�		g����#Cz�i�mőO�ǢQ��x݂�E?mŕ��}~��×Īt��kC?z���IQ�wyw��?����%6E.��%_������ޥ��֯_C�:�R�46*]8YZ[���w|b"ɩJ ̝(���$]�}�wAXɸ�i�Љ��\��y�*5�GQ�v'�<(h-MB���F�B�W�rnp� �({�dl�e�7�����1fU�I"���/)()��>y>��2�_�lW�_��@�Q�F���7��m{{^-�Q@��::0�D�+��_?����k'w�S�o��z���x@�~wljjr�ݜ�1'�8������j��e����ʊ<V��z�<30W�#�$���h�޺Ep�A��������k�bw� 2���R\��\��R�]�O�A{{Mv9�׬I�s2������;� �g�
rI��^�ss3��$s����˜��/W9N�ee@�O�� ��[�2M��g]>�������d�QC��[?@^Lݲ�2_�`3��p�����^�/n<_�FqA�m�㆗>o�"�Q9����%W ��Q�^^��i.��k�	!!'^�d.�v����Fұ��NMMES�CK�SO-嫟�UwX���!�s~�/�h�J�1�F	ǟ����U���ϽwV�iu�:��S��[�;�"")9訿�W �H�͚��:�y�&[1ݩsll3��^:���CM�e��]]�+����w�n�.!#�
����K���Q��~��e=8��h��C*�b�֞"A,�Q
����e6����+KKKlŹ=*��cЉ\^�z�r{\V��gf�<|x'������꯮�pρ��=��7*>���gj�}�����G�˾���Y]�!��^��w�w�!���ӣ�I�S�pop�iFRX;_���MWJ��a�2���
<������³�:ϧ���F�������L2u�������u%%\���/�fh,���?2}qppx��&�n�S_��h��SY�sk��0T�L��A�Ȥ�����*�;��ME.?Z�7,q�>�hFs�s@n�&�u���Wc�IMz)���e@���L8��	�3����j�dK_�	­�����@2�#��%=yr&Jb|������۫c5|Pj��'GY[<+�S/f���7�3�4{L��6�N<��z����,+^�Ko���ё_�����Q� re}�����0!��:ϋ��D���@�y���-�NN~~�ci_�_�uU�ΐ�د�l���nn+1f��J���>[�ܖ��,s���F�ߕ�o��{�4�Pk���bV� 99��c��3����m,45)'��'����A�;���󜜜�Y�����_��6���y�;�e��n/�{�ˁk����y��4s�����a�A�,ZM��n���[��T]·Ƅ�D�
�@r�*�����|ƲY�9���8L[�����ŉj1�%l�Y}֭�?_��/��ng��]�����$�;��1w��᫭s[��������yȚ�(�th�8Ă������������Z\�ZB$�������[y���W=;�$�P�L�T� �liyy�����' qk��ш�ẵ��L\�,AV\��LN`����wK�@P���.�J�O�v�.�ꢹKK���;]�T�H�pC�lbr�ܣ����A�ҶcU],O�8�����M����A`�{GPMῄ˗/�����v5�rY��홗*�躙�3?��`�k��=��Q�4�Rk�Ŧ���\�jH�,�J&T|_W'����p��*���w�޽��u�I������`\����_-Ńe"�W�a^vy��3�0�� �D��"���F��-��5�_���))�Ct&UE���!�T�W�HSsȿ�e������ɓ�-�o����a�����_��6�611���4yH��P!�/Z��������=��&�د4��ś_Y��Y�%��A��&w����ݕ��_�����T���V	z��拊|���@��sl3�C ܳ�I-f%��1�!������w֜}�	��Wz��֠���<04|��bv� ��
������k	y�.����}��U���%Pѩ�1�7s��;�����*苫����˝&�� ��������",F�a=��x���!B�Y�E��_����_x��e��v�/��^l�z�l=8Ftim-	��-�����/q8H8�1aII~H���ޏ�n�Ծ����w�S����FHfKvQ�(d�̲�h��X��!$d��8!d�c��� !J8v��w�ޟ��?=�s���^�9��>���6��{��δ8�:$@��G��o�l[�C�8�W~ծ�U�.�2�l<�R[{����T	�yX�����67@�@Y:::��p[�Zj#��6~JP�r�&&J4A�L��y߳ ՚�(yT�[�kF1ryp�UP���g�[+��nP�~�%@����v����绅�m���t���m���p��h����M^0E�Ü1�j**��`��?��x5����۟���"逽�N�!�w$%y�\�m����gAk�_Q =-�)�[���k�\�ZVޛ)�o%U
�>`0.��=���򧠠� t}3�7ۯ90�M�g��}���T�^~�(��`Feo���Q�ci;n����f�v�8��(��O���&8���^*~6'�F_��* �vJ~���7�z�� �/PL��Ê��Pz^��LK����urdW|���h�xSԛ"ͭ<C�w&�`c�xM�ΝDDD 'E=̍�-[Y|绺�{	�O�-�P,��+��Uy). � .&i�S���~׌�Y{�X��]��ln�115Ս�u�����Հ�@$WGoW�)P�����@&dX����i9�%��oӨ
��Ԃ����GF�H�R��S�����M��Ӗ�V�>7��H��O����?@6xqۯY��E�uss3\�^ a��Kj�s�0&V�H�юͦ6]oڼ8w���i��*|&��K+��ՌNL�M'>^#88�L�y			|s
3+555�X�b�ȰM h�R_�2�$�I�He�}�p�~BV����M���U�;��@�}S����`7*7[8	\VYy�f.0i�3�6����q"�.�~;�&j�a�?�$\k�9�<�.�,;Z)$?E��"�ִWUc��嬚۝&H����|K�u��p�yQ0���k�Tuq�����Ox{����d낍�ֽ�	�l�Io?'�WT9�)3��h#� ��r�`�
��[[5���=�t{�թ��٪�5�l�B.Ϻ�%�W�4$�ӯ!��� 	�Rc�0R$����EL6�U�5�3�����dz��ѣG0C��� �{�U,��7��Y7����Ћ��D�4�[�{�2�譳�=P{\���w���K����2C@@\RRR7�)�?e�<�v��h��lAM�z,9%%%nD"���`�W����,[�#.���8U�0`P�l��
���U���� W���c��g�_�<�h��S���/ook;��Ϯ�uZ�:X��G�QO�� kĆ)��0���-�=�2.���&%�a���G{��o��p����������N`���D6��HQ:��l@�:�����z�:e�=�A�0���7������yM��?��J�Xĳ�J�9 u"��	
��%��fZj`V��_:�J3wf/lؓ��A�M��^�y
�m���I�5$�؃P����W�N�a�Y3r!�.��0cVVW�~�z�n&����r̷6�xUUU8���pf�If�k�U�,����o:��6$�NNNē�"���j?~�1���|��=�l��/�<Y��=*Tx�l������|m���C��xS^J���/"�\�;��7�G(N��o��cggG�������- M/��rop�5��9����r��%|��I%�<+ӫ�E�	~�����	`d�����_��wfgR��O����!cE�7a��\����tڔ��ǗVꦨ<�~�d��askWAGo� �VS�lΤ���TOT>�c���Z���� ��@7��ѿ;l�����
��?��d�76̪i�n�~L�^�Bc[��1�[����SSS�
�{<A��]_F���&a%Bl��=[���ՠ��ԮuPP�uf��&�vx/a)n��"��"�x��a�]������@|�H�Ȓ��%}�wg9��ٙ����	z�҄Rn�kk� �	�m %�����[Jm�W[���ٹ���>f��,��� �k+���@��<��bSw�9�V�Hv��l���E3�`������N�5��L���[������+���h���J��v��_+T�G^���eN��p�����P���"��+`Sj� a�="��W�Ԫ���͖r��[�P7�:,��Uaz���F0�e~D�~��^��j�W��K�Ė*��п��/��h0��N����� �.Ԇ!���mnn�eeRx����L��|˿y1��6�hV<�h,��_qx�zz��=����r��Ƴ��
:i�-�7�E�?~$�Z �GIEE��('-��d�̇���͉?/��XN W���챱�6"�m��9{_9{cl��5=����s��VB�����}��|������t��k��W{㣣���'���Dl�1�߽ �۟�O��
�n������`��2;2ΰ�?����y�_JW�ϩ)�kos޾A	�v��E X��;�;��� ��?3�����/�$8��^���d��7��+�����(/Wo03��#r��d?�h���"Ӳ�/�Ե��C�r�&��\of�2j�WHJ��� B)��$�s^g���pE�ݭ�㆜C	G���tp�Ys_�p��B �%��`����I�ִ�ފ1PfdeQ�9A����V��R�$�|#�Cs�b�~�s��h�r���Ӄ
v_\?(<CD�m`)i���@�w�����5m�GJ򃁓��|�6+���Msء�fX��=Kg�s��:@��F������ xIZ̿�<trq����R22��;��W�Zx
�7q�q6 ���}����::����924ϜK�ŧn���1ZO螵��Q�/���^^�������t�,�^~&s��G�`�c2�$%:s��]��UV^Z���lR���<eX ަ	�WU5W�Œ:�L�rr@j��jB ���TX�EDD�]_��3��fE�C�q<�`�o�GY ������E�6��+u�6���݁���Z�m����	�bN�E�P�.�;.���v֣P頣����Wi/�f+4�D�/7o�Z_���>�Å W��l*J'�$V�b�p�0ο�� ��[s�
��b}}cxW~����H9��Ӯ���G��'� =oo��R?KeOKM%��+,{����Ž��FP
Etx�CYY���*QP��/`�~�T���`�C�jС�0�
&�;�Z�t�_u]�ԵvԷ���k��f�ɬ`��"��^�Yjo�,�*Eί߽s��~�x�Դ�{oi�6���$��bbb��Bv c�e�K�'�l�{x7���~Ω��4��5��Z�f�4��F �ollmk��7�G�<����S����������c��
���g_^&?7[��ק"�-ݯG��X�hP-N� ��:��a�;�k�Og�����ߎ�M�����--�g�K�X��1�ҐAX䛗/��Z<���\���Ѷc�W@�9��J!6�'��G������R�I�` 7Mb������+<f��vBL����L�aE%����
Bəb.<:����V�e�W{�b�=Un/u��邋�q��w
���?77��M"�@��4�Ʌ�ů�E<��c�c ���ｽ���9���$_8t�5��T���ĩ������$�?r��H�W�9�d���SْN���閛5Ύ�]��GsZ�������������	�Ȕ1y��唹x��Б�D<���C��N��A��,5�-�j�u�o	E�**W��]{
�����6I�Pp	'�,:هAm|u��Ç� �h}�5�II�w� �<�T�9(((�Xj=YJhnQGp��zh��6�t��Ф�֋����g[<)/���#��!y3 8�3��O,.�d����U�������;z��4�u?�;�vJl�Nm�����ӧ��`W�K6䇳��me�*a���� 6a���)d�����Ibqsu�I���H��'? 7B�}��ϊ�4L�T�TIZd�aia���e_�0CXxh����L�j�B���QZs^�[�~�qC���r?B]`p�t#kc�~�
:^�<Eט���`ychdThXʍ����\C��3, �3�߾�����KKI�F<�RP�wR�L��Q|~�Ҿ7õ����*Hh�L ��Μ�����*�-W7�?2�-�;h��_���T��zF�A#�4{�vd�v���F�`��A���g���D�3�S$��Hp�R��z���7��o ����=10@;���,9�86�Z]E�	+&����б����Mh	�4N�� I%sS%�v?`j�/[G[��W4ʔ#�<�'��䫄��SFFF��P1S�Ǐ��2�^z�H��1��um;;� ]�JF�a|��n�x���,5`3s����Meiiɔ�!)	�+��t9P����0w�) 4p:���#�
F������K�T���+g(���O��������A5�D!/
��ȟ�S]�u�XN�F�����ݻóc����B��kk� ������B�.7��	�Z-r-h��Bb��S6��p��!�� �M����@!��6���G�<�,���:� ��_��'�抖��A�)���G8E=A�N��4�{җs��UL����- �j��"���}�ܬ�g��:�����D����y(������$����̎z���~����O)߼�}S�{��z��!V%]0Z�hs�i`�+�)��D)6y��]�nja,
�L�F����������k�SS�Ҟ\Y�i &�� ʗeӔ���g+�'����SW_��n\�ʺ�ݻW�/~jh�l���Ҟ^�q���t¼l���-Py��@���O��1���>Tbs>e51�;������/�L��9��/^�PL���w������x{�:��0��lo{�����8!���ɱ�e�p���G���J�@�,�%ܪ���0-34����L�޹�ސx'E���_jWZ@;�b�Z��9|�1�xk�(����h&P�O6-?}�D�y�,6ut��ݟ~z����_Մs����ڸ�0o����ԮmTnv�	�	oa"�!(�?�����td�
���+�����6��iC|Q�S���b-��"JJ�|lr��1�s�VV:�j����v(�S��A�U|<�Q����@���YwQ11��!���kތ�����}�+&�6�wc��_��C�zm��/�xtT�a
�W4�E>��vv֒��4�ge�~�B{��4A�I��IzUTB�����/�6����+	��h�/���U�#�Vl/���#�eK�����' %���v���a�S��'���'3��%Ϙ�����&H��S)���·��c�C�{�}�7^ҭ���44ܟ�}*���ښJUQ����i---q#�;;V��R_�	 WY�M9{�y��XZ���,A��=����r4+�*���:[kb�%����m~C.�O--�)��WcL1�������;;�]R��  ���CCC� �{���]�cKx�����b�"�Ԕd���x,٩kŭ���b{�-���na�Q&L�x�r6A���PH*�@��U�l>>��j/oęUg*X���Ǜ]�uS0��qc213[�Ә������n�Y��2�����+�����!(�D��sz:�}���<''' %����rE@� }ZZ���P'o%UZ΋_�c�k����o��|�`�J/	�9�~�z���_ K5긴��BӲ`�o��֧��l���2'��?����M�T[bz0�i���D�xi��C(�3)d�,p��f�?�׫�����=���g�(�[��>z�S�2�ae,���IPs��m�&
��������2����er�
V&&.�\B�qX^��1]n�PcN< n~,�['�k'��5����_�����'�T P����#�>i�a����W�@���08>25���A��V;d$&�s�IxTxb�iH���QQ�w0�_�Q�ˋ�XXXh{	?h����>=�׮�Z �Gc}������vP�G�W����6\>���F{��k�6}�S�C��@�~���5��k���PLu D���7zȞ Q�^l�I0����:��s(f��s�����0����|t��������R��ɖ�S��
�0#g��gP��>֡^�XW��kS=���Q0��:����G.x`}>���(�n''���Z�q���w�wc�;Q%e159�
ڊƖ��?88���R�(7-s�]��õݱ�5  �@,�ák<f�cɕ�c���x�!����6q�1��'�=���gjurw�M�|�>qp i[��*�i������~�vd"�+gm��x��8emK�@��=�rc>u�LJ��_����Z����PH�k��V��y��ٰ�I1�b�v��{�⇞�@MT@}�����[ls��.��,���#m�'�{�꽈��-��u�����B�eO$��t�rS�����%���r��5PC���s�O51�m"/����7���[���D^Ŝ�mlE��@�B�^�A����N�nh�{f���=�K�B�0YY�_ ?]ٜu5 ��FGɞ��E�1��`���J�?�Z����?l$5<�sm�~T�̢�(��e��A2� ��.�]]�ͦO�۸�>z$\�fV�Mw)w7��ԭJ

,� GQQ��m ��c!�$m�[���c��{�Y����<�;g�o���A�ׂO��(�)��m\��4�#�e-v�G������4�$Z��AQՠ��V2����E�III��,����������������2�9%�~:c��{�hg�U@]��!�B�%/��'E�fG�ONZ<� 5�d��]B�o�k��i����7� _~QN����/����I�����P�����ӣ���D3C9%��]�=v��}B�_Gw�f/tLS$r�����4"�t�A�a�.9�{h'��pi$})���)H�XDZ��ZH_C�|��^��[?~|=�>/S�����Z$�F���˄�u5Yo�vT��у.6 }0����ɥ��7�&��I����.�"���"&�'Jl7���J�B��&��c157��R��6�/�U��ׯ_Bei�*JA�l���[��: �j��N"ZA��s$1W���^�B�3mRҔ��m��՞Br��~ ��&���?攟���s�m!o�S� ~K�4�n�{��n��HY�iik;d�נ��l��̬���+> ���rz��GT:��;y{U��=�o��f�|l���9��O����ަ�#� ��!�2���pQts����1�������U�Q�O�.��>I����H��'�ַލA������e��"�46ሁ�؅!�lx?~12��8C���bAT�����q	+��9y����N�W��@�Xs���	�T���t��J)ƺ��g�������>���W�Ƒ�!�o`�G��g�.ːB�L�}k���*��?�X����EYԋ�n[~��1۰�h�.7PmX�@4u��=z$-A�T���C8D	$��=��-��"�'l'�F5nMo|�>���q%�(���󥄠yT�����cA���m��5q3j S�T�n���ff�m�Q��򝹘W��BB�����Q��N6�
����o���o�(�-5�77��E�V�m�ԋ	�Aí'��2޵�?a�}qv���IDR�,�q�=�D��g�=�	���p�IT#�1���x �Pӆ�G��}���?S}�QL#SS��VB�e��%��A��'��!0��b����v"�֫"�E�76����^I0�����m�?�>�M<�A��~�,'%��LM�v"ۦ���Σk_�}l�ѹy*���7�6��&'2 T��}_Z����.Q�&1�&uZ������Z�:�Sp)w���u���9�����ř��[Jl
��_���_W��MJi4��JoDp܅ �&��`d�|�mZ�\s�P/Nӥ��^�`�ڟ���Bd�xoA�SqJjj�*qI����h��Yw�۷s��*Fjy�d�70�d]����U��mCx�8�<�YXԯ_������*�w�����B�O�e����a -Sޣ�ޜ�4���:���Eg�.>@��߶�����e�p�F�� `uM��H��FRV6մ��:z	�$�<�"�[�&�v,�������/��vA ^���%��]��#{B� C�S`�?gH�ڟgsߗ>���.yn ҅
��P̛نwo�@��),��;]��z���b�T]���#Ҁ���I�]:��c����(�=�����}~�:�_��f>"��J�̍�o}G89!}E�/

؁�;��L�!|�W�ey���5љ�H�NϮX?�8"h���"@�@��A/��WVV�@ �_C���~�����в�����3���4 ��������l�Hqo�v��8��>)�o�����W��1:�g�}Ey%Y����7�P6�VO(�Dj��q�ߞ�	���&���˗�gv�D���ֶ���g��qpp�}zU��L2���ͦ�6��-m�G(��~�����~��A���`~6K��`�"(k�������su �Ն��]�<)���`����p���v�ov����a��1� lf0�1�T���Ǫ����o=:���Xm������`/�}�1�:��J��$	kck�������?A��ihG)=��L-k�r1�I	'''q#�S�/�!��/^�LP�¬��e�z�@���o������^W)�7�i�WH_�wZ�n�H�����ꌉZ����x�0Ѻ��Q�g������G�_	H�J��#�:Z���I�5�%���"mռ�ĳ���Qو�C S�S�ӕ='�L�>�=(<���X��j�Oqt�8J��\j����·�	p����;��
\$@�K��V�d�	K�S�#������v�>��F7��!)"��������O�]I�G�o2�0�8vN���ǵ{��u���쟋dsl]^Y�wS���p��v��S33:Vknm��#�{?���1#��i�>ϜaƉ.Ԕ��'��s~UՄ�-1�A��t+A�n�H����mR�ĊnY��L������i�	vF�J���/�G��N�x��mф�Qv�)?ȱܸ۪�i_�ܛǸ�#2@����.�@�� Y����	[�������t�a�m홨��%��a�μ����!�T��9W�	E^E�P.J"���Mf���ꕊ	(9���� �a�=��ZW�����n��=`���hDչ�Ǭhs�� ����$�b�����r ����ف��� h�k��� ,I��3"����*BC|��:�^;O~���]��e��5��Tk�e�}������f�0�.�S.A�uIt���nxS�V�_w�������.'�I*��H���	�%$�DHuў���pa?|f�VR4Y���B�A�~uc��19�2~7���y�ߺ��!m��L����*x#�����EIz���ʊ}l��9yDt��i>`�R+�55x�=o/7�NQ"��fΕi��cx��~��Hp�C-������b����]�P�p`s�a��h$"������������\����pH��]w)�DS�o��g���1��J=��-~g0������+�-��\���U���	�^;yG3uS/�D���<'!zi|^sr��DG6'�J��9-�Өu��7�.d(��w:}��+'�Q���hiF��(��i0���+-Eu.����k��i����0I%q�����v������y`=p�f���ڱ�M�k��v��y��s)zG�@8��� ��M}�������ئ�͵�MրS������$Y���wD>�M%""
�]^uu�������X�YaW���c��d�`&p��(���omPV�e���l���O>F��nxQ�h��x��p�j �x��*v �9��ĳFH'�vFw0f	xQ`�:of�Q*����q�+�,����g��i³{�v��ETQkӃ.]j�85@]`fw����p>��ۏ��!��m#��!��l��	^���w/����P7)�q�衈8Z�R�9loni��	����F ͫ����hSX����7U�A+lB�O��]��E	����"� [�	$w���x�Z���BK��Z@Q��IF���a�>Ԫ�e��eP<Q�1s�w8{��Ĥd���a���2 ����/��%���gQ=�����b�N���lC(��a�L|I�c�n�M5����՗kd�Sp�����'��J�e���������f��0Y�u�8ez`BZBC	��&NW
����())#�������?�,�	$R��jnԐ�Y��?3|~X��ۘ���Ӟ}�b�;��"\`I�ǚ�H��(�kL�g����m8�ҒG(>�y�R�ǗIA;�/:v
�oV�Xb[��S8��M�ꗄ�i{���� ���dw7��JH$�:��Jֆ(�z�ЮPC]A
V������~����(�M�忁�Gz@�=���q�˥.r�Dk����XP�&��'���p�W5�<fl«}�ã&��������Hg���Z/HBк0в��;��Ɗ��)>]L_����Ym=N;�Y!�h>"]�̚��w�9$c�?��P�E���>`K��Yl��ou��:�H͓�ֽ
���æ��&Ay�$S� ���n-că?R�]/D�x"��d�-��wt�	&���R�E#[������= ��nƖ�[�sK_����������b�<Lq�:�t��i�����L��K+S5�o-_���N�X����P�'�Q�9���j����k���� ��	�5t;�a�ɴL�`��$������}Qի++�<��ba3��T����t�!�����2�B�-dG�y�2�����N���X�~���+c��v�=CA,L��[��'6Wv���h$� @#7�iG�:b�N#(С��zA�Ǒ�4eVB�����C%)))�p�NN!�` ��e�6���[���l�j�ު�4~PRҕ7`�z$���u{�����f� h�.[��Ha�����=�����wzr�4A��]��j�
'�M���^媘J��Y�yǻ/w�@��ybF٠�;9��^]���/�@~�*{�9I[,X:���C�&�
%���Kjd�����	�:I�%�����:�'tZ%_�$ƃKƙ	��7�-*2�D.+�3-#��l��K7՛2�]_��).���[������ ��ldX��#5.����b�Fhe�PcM~G[�&j4�~vc��h�!�P���$C
���E��~]�,�!��+\���x�9��� \����m�S�-!��	n���tP{�'��W�g:��/�~�lտȢ�џ>�����:r3��A�U��k$�N+]&L����a�{R'W�kzx�/�ί�5ľ������Q¯���5qʫn�w�V�|�H��1K�_��|s�:��Y���Ռ­r��
��Ub�\A3!�����mt�^�V�����
��ca-ٍ��A~i��L�}�[�_MlnK�{+�M$�G x���d��Ӄ�q��^}9TV��D��:���4�;˫ �/�B�԰���@��=��Ma�D[�<-k޾�>Wzm���h3<oZ|�P� Þ��G�:��#d����v��6k깾��i�7{G�-���(���A����$�$�����-�^�{O<�-��I�l� ѪeZQ _.��<8�O���Sq�[��y��{��xd��m���Uҩ��pp��GTcg� e�0��M�<v�ώ���_����o�����M���/��T����m�ڷ�R���W�/?���|!�_�(��d�;9x|���\�<Pd�&s7C�-��H�#}�J�k�[�6��!�=R7c�\��P���4����E+,e�aA��M�V
�)%�?(�_�j��\z٘0���ȰZ4G,�=W.�#��z�K�X?���Q!z��~?@֒y�D���@ˆ�+��2��673�PV9�C��ـ��t?^hw�@r����/2l/�/���t4�V��^/��Ѓu�ǹ&P����x'��9%c1�����t��3�Sϱ�!H��(]c�#���qeR�g�<��Y}�fQ��(Z5ΩOP*$��`}��S�D\��΄y�)oK��8n��ɗx�U���zP�\,Sk�Q�Bh�K�#@���m�hLr���Ō����m�*���K�U���vN�ϟP����nï	�z�nzS�o}�ӯe�q-⺼X���k䓁����ߔl&�f��c/�J8֚�9l�iL��.F|� �� ;��)Ϲ�ҢT���K����ǳs$��B-y��j�`�W�K���g��ֲ������	 yb������D灡2�8�v�+�~h�O�u��2xx�\n��W�� ���2n�!da�r5�:+�l[dH6G�lW��1Px� W��AJ����u�~�J�Ǆ��\u���t%N�U����)��U,�/ lZ�'���*P��e�uҵ~˻����i	a�=��:�Z�z�
��&}��bt���\L��B1}Piѫ,Nl
TC�)�r���b���|s*a�E
^�n�����٩]-�0!�
�ަ�+ ��i�J��c��������"o�-+�}�p�����׳��nΟ��* ��p��"Ck;��5�6ĴJt�P2y�B;o)��)�֋����@�k#����*� b�G�؈���`�N8Y��u��lJ_�&D���J�V ����÷�T���B�_ߴO�%`8����Ǟ�	���}��JR��]g���U���.'��ae�]����wv��Hp�j��-�����T$a&�o�����/��p��J�@tmb^y1n���('�Z┞�Ft�^�[
Iׇ0)o��l���י��tФJ�����s���1��9�~�}bD���>��O��y_��kX7J����x�@LΛN!�|悦��$�]cH�[%�Y�{ڀ�)tEH��������W"��(#�<\ΏQ+l&ts�{��AZn?K���<�y��p�t-=�ҿ{��L��?�b"N|8��o蟽+�'���,v&;��:�1=��a��j�v�_R@\'�?�R�����IdX��/4�Q^���/�n����M+�'�����ڳ�����.��8�8�갆������h��M�E�רyK@�$�ލ�.]��O;�J�'���&�H��KS(#\��ua3����pީ��R@)S�+�𓆉���;�/�������N.���2��ꘅ�a�1��A�ܳ���s<� �ƎPX�T������a�&ǽ7�!�c�]cr�%�e����Ǿ��n�V�����e����\v�Y�2�4,h�C[,�[<�<����^&��%ed�p��b)�c�ۿ���$�M��g�!}w9��y����"�I�簼�����'������0�������F��$@p��Q������s2�9���lK�q&�~ډ�|_gz"+������Fr}f($#�/6��d�u���%=�2~s��@ZZt=��.��0��{l�,��
(&����v��K��������-?^��7T��MK ��"	��VퟦZ�'Bv��ݬ��j���f��OIlYӣt�F�J��^�P0�^�.9wY}�b �D��_�];��&��D�~�cX:LXa+���L��a�H����NL�6����R|�i��.�Q1� H,Z��A��im�ҀQ@�+e����5�Ak�0:	e�{��(�Z!��T�;f�D�1�����J:`L�+v"]//���G�#�����'V�۵3
�p� �Rw���ղY{TC@Mm9ӪO���ݸ���;`6&
ނ*I�	(\P�g����p�� ���_�36�r��|���B�{m���v�$k�ts�����m�"������5��3�T�5f#.�.����h ���}�,A��m�L|&Ͼ��m�#�E�ߍI/^Z F�^p|�������*PC�I@�ȫI�?���ċD�1����;!5
/h�L螭��v=������H� @&�~�.�*�v�yJ�{z���&& ��!�*!ٝ<0�+]�3�R8o�XЁ�g��b� [/���)qvs��|X#3�3' �>q	��M����$e�7O˛�f~�z�Kƍ��M^¥�`�:��, ��"��9�/�c�!�K��z�ؾ�.:~*��¯��'e�]@Фg����`�r��X-�r�:y����/n+1���#����W'����'���FF牢�]!�>�������%��Oų�`b�1�g�,l8��bC���=�g�O� �Ն�=�[��/����83��'�Y;�]��	�?� P����Z_w��D��(0���aN��hGv��VG���	!�Xpd	���B������M�eB&�Dߜק�	T��imb��l���:7$���k�<I�tA��+W43(�冎��1���V�o紸�v��) �h~o��Qǝ#)�jpT�z�<!R�f�w|���������hh�_��׀�&�����`#�t�z(KIA���O��G�7�3��;����)����8��*=w���kmT�FFG>�����{���J��ې�����qʣzp������� Y�q���y�_�[�y�ٱi��vKRt�9(�G�A����ݗL�ðU�H0�w�-N���Y�T�R�ϕ�^f��`س��0��VD����-���f��@P����d����*o���6��$@'��PH��3�#����/Y��q�j�#a�J]Tь����݇=Y��k���R|kJ�I� J�)����G&��T\V�j�1��*�Y��1C싟ՙKh �� ��3�s��h:�+��R-O�v�B���K�ϡ��b�py��h��<99�����}|��-���sΎƖ:�Q����w=C�{8Y�[�=��ۯ����P檱�g��wU+�/�MS��Xo�a;e,`^A�>~�,�2��7e{6Ѳ��E � $�SJ��k|��
d�
���7���py��[�*�g�x ���H�)�~"ل��gd�����h0� �쏽��V��O�`�7��C-�M��rʘ��N��P�	�~�u{�V�.&��N_C���.��2�ٜm��Q����"�j�1u��a�P�>����%=��ߟ-�.�)�
k�N���e<��/ϛoq�ԩ
Y/onv����܎\�$��5��M��]	qq�"���)�!c��qJ�q�߳I��PĠ�s5Hd��M��V^�i[��՗�# 2�Q$	�� =@��P/̯���&��di"� �ʁ����!�wCm��-k�N����oe59yo=�����m���Udd�_�R������@ɨ;�Ku{��ve� �Ɠ��'k'E�O�J��Y́�h��U��s5�מ�5�b*_zs�<H���ͼW��������g�=��q��B]`�c�K��eF��~`���nO'i���MD�w�񃈈�t���t�P�
��<a�UCL�uq}������$6Xʟ�ے����Bm���p�︺�Ҍ��=�R�t^�5i��ԉ���VD@�7����Oa�/�PTp�3A�/���Z�z��:|8�"'y�_�$�*PA��<��x�����Cl���r87����y�;�B�(���7��;#���y!�����L��gq�-Q�i����0&B���a|��t᯾�ߏ'Y�f�vE.��`O�O�A���CmL�7>�+?*&w�%��H��h�2�(}�,�L�.=a[:�Z�ٳm���|lKY^G����
��,r%}偁����*.y��-�V�}mD%��Wg�x{��#�`�$��xS��<��ͮj\�b�U�z�S�犛A���s�$�����!���wد|�@�U�FF���aʷϳ3�Y:�,����U&�x�s$�����|Wk�4��<�|�<���9Xa�j�[12�'!��f��DiK(CsZ8c�P:��y�T}��<��qJlyͪс�x����p� �����u��ܡ�4��ܼ�-�wC*�n�����K=+��α���	��Ը�����~b������U_3���G��:q�p&��yq�u�^xj�j�	�� 4��t��k<����J���u��l���˗�d�1�X���:���-�hgC������U󝒒�=�����y8*�r�޿&��࢏��*+�ɞ�fi&f��Z՚6�X�w��Pv��i�<�}����3�� �HL�g���1avO#��T:D����S���j�z��'���N�v���y��y��4�i�wɽ���:w��W��jx�a��8�-S^ib螎��ꉟ])����]:��t�q�h=�3s�J�&�_uIY�l"����J%���y謭�����x�፬�T�����]�\]�nq��z�K�6�UaΈ��KH��"te�}N�m����M�hi"�W&YbUz�U�k��yQ�p���͋#{�'��$�����Z�/�a�,���a�C1~��	�6t��Đlll�	����%M"q#����B�X-��:�ID�z������]o�;����ş����ez� ��D
���h��gZ�SWR�R���v��gV�|����6?>��Fߓ� �;�H�>�9=
Ɯ8�:� 	�J��s����դJn2���{Ϛ{���,s5�R⢟S�?��l3�x���H�3����s���V�1h�^Ps|�ǌ\�u)�ʖ@�DG�������TW�:wG�.ա�����#����k�GZ�M��_�$�e�r]~���d	 �!��f#ΰ����pj":*JSie�OG��1�QǨ����Yb-�������߈�hR��j."���Q�����ig
b���7)�͛A�`u�_6v
�w�f�Ϲ{z�Og�b:r�fn����XU�Jc�嶵m?�KYQQ� ���;�4��,��j����غ�;�����;�B�_�LJ=���Q�̈+1ʓc��LR:�.����X:��shh�)������9�m"iڨn���?��Qs2C��/4�!��˻q<�iı���h�+īHcT@�su1�hmb�'��s�Q���Cve� ��l����v �'�t%]}���=g�.�`׽�p Ժ��m���z#˨�F�M噕v��u�Ҙ^UGeɤ;�9E^�T�%�̑�O�����5�B�<_�����9�����7a��ݨ�[������(��Hq�����.�f�4-�"�<�-��&m<��O�%�Ų��grn!Y}5T쓜|��GU�%X2�lmzK���Ne��'ÞU|t���}�==���i�G���Zړu�r3x���F�zL���MIf��`��P��O2�4PC/]�5b�E�x��LӜt����ܽ[xOik�x!��̿�cw�z�j���Җ6���P?���V�;'ޜ�l4���ek%��&W��>d[b�W4z�m�}��ow5���jDtT�w/����,�an��z�Ed��Z��~�?��%4�|n��J��	
�--�����G�w�c���K2
YIVzI�����+�=3�{��약?�"�������C2�����w]��է���x�����9+����k�?`�p3ɝ��Y��힣�c�˒����\�-��O�Zp��,�$G����Zfh�5r�����HIW�c&6
K���������	�q��kU;�~��^���Hr����CϜ��V����m^S=rt�����=7�Ru&(���k��6Ӟ^�O3$�%��F�0�4#}�l'�����������^�]eפ.Q��8�x�ډ��$�f�
������CA��,O�ĝ-kSvI�#��GGz�z)�����TƼ^D�xnK]�8�������������"���qs39%�Ɖ��⓷���k�9 !dӖ�$�u=����<ė��b���&�6G���,|��h��TB��۵��Y��PK�o_&�/&?�5V���\��I�$�ux�W$jh��(4TU�\���^�����b�.BYZz�o�f�O�$��ö��L�aS��s�B�n?˳�{5;c��6Z���̫��6wsy��S��6M K�|�Cڶ�D��ǥy��ͣi�T�F���h��UM� <�	����Y�A0�ҳ#����N�s�|�"��C2�n
𒾿�7
��MkPi/�:�6%>qw��s��x>�~����\��e�����qIP��a�I~*��U�<L6�]����޼�(���җف_;��h1|��ʘ��$OƝ9��A0��/�S�@�`E�n.����ť�U�i����W<�º�uſ�j&3��(���,J?Z-/���}|Q�@�������'�-�~�D�zu��r��w��i2,�"��g�g^0|\�ٙ����u ��z%�y Z(�xx�J�[0�މ}�wz��O�|t�T�l^�� ��xS��*��k�5Sn�)L�AE,ն����qS2�Te��<�i���X���`�sV<�K�1�z&n�o�#�3;lꯣ��kޞ�?_���.�F�vw�.@1���?��NuP��E%%�N>���5�h�[(T=�fZL�#�,�T�÷Gn����Kť�F/����:��?����o]s��~���������9��)���_u�����\�q�|>�Eh��u\L@W���͍���m?;��W3h�{�d���dd��ߊ��q�C�M�����T��vcю��h�^su�2�����<ʥ}�Y��-^6�<�(��P�;�!���v��fVJL����j@�\q��
h}�F|���E4r�X׏Ҳ2�^h���u��oMueYs&��q6]�h�qR��;��*�R����ˣHIG�Pd��`x�9��j���Ɖ� �W��m��m*&��},�BAmF�q�i�9�3��'''YK����P��{��l|�������W�����Fͮ�6����gg���������2(F���~YZ�!5�e�D6��\�҈�� ��Xդ����;t�,���:�K���̱�����w��Ym������1��q�D.�X�Ֆ��L9GT���$�s�4sݿ´���vpj̼��u뀑Jc�a̮�o��ٹǔ;<U�a�+k
*�Q��B�#I���e�UR�a@^�f�0�Z&�9	�ZT/��?��W�lO���N'~�ǧ��lɍ�ss(@���ƛ�}�����]/4Ny�T}�x��-K�- �X2�|�X�T��·<�b�̖�?�@/��l�EC�]AD��h�#iu3TrJ۬ʉ�Cc�g)�/ڊs�G�#x����L�A�C����;=e�m�M{������%%�^���K$��.��)���UaI���CS�Z�Q�8d��C]_45E�(ζ�������bQc�>5�ݷ���J~����3�>k2�c����𘲫5�`(�_�.,�4����[6|ssި�ۻ&΂k�C�Be[u�>m�gyIl�J���[5����^
E6�(����ZE�+7Hä�v��~%��H:��ɏ�ƥ�r�-�A�o�<\\���!L˜��Z�B'l[Yu/�T��ΐ��g�E��sL�>p��^{�ǖ���~h�e����5[���N�Ԩ��s�'5zf�6�O��q�ѣ�h����W��(窉���
(��.���bej�YQs��F��CC���F~c����N�Jq�����x	�a�i���Y8��D�w��wKg?P�P�qLV�m�݃��!�,����y�+�D���z�X�g���w���hm��s��3��{�cF��7*F5�9謠����-y�(T�fiM�M9;O��q�T�q3��w����vc.��9�\2���WWڿ$�T�%[��68���$��X6*�]�$�~th������h��C��/��N��*�ͬ�h�� ���2���$!�fP˘��5@'�]�@��׻�[���k	Y���]j!!��&�W��/�j.�GR��0k�U*��y�W�4�n����7i	m)P���/)+����ZTz��]�蝫/&&���揬��j�*����5���ݻZ�%�Dc�}G�N�LWg��>�'�����q���e�)oh�Kt��h@���:6L�v���B��U`"ϖ�0�����/3�����L����#��e��~&�+wG�^�ںf���ә�0iWk�7Y!��g��)����6~�T���UP��zv�\��to�6�.��\��G��>>F��}3y��ϫ����.���O��̑�Ğ#/wI^�Kÿ�e���)\�.I���]�}"H���������'<w�T�:!c�)�wVq3��I`��N�j�_B�lE�5�7k�n��t�6�"zB\����D��?�z}%qH[���{=ܻ��S���:繄	���:�S�q|�l�BD�y-�h�z�8�h}ɥ��p"U@���A���%#�V�E��,M��sR:�,�Tf�C^$�1���7���3�������s����&�[�8xy�m׳���pA�fu�`0y+U˿s�+�PI���o�:��O|����{)���ib�xwb��%�#u�ZL���V&*2g�]��4֞����~i5�͛�)�pi�� ��20����u����sZ���tY$A�f�)*��A#ܒ��Qo���~6 R�|-���xĥ���@�m[l�����2��\�ao�ی�-!7��C2�Bۍ��׾,p�'�:K�~]��OOJ���w�~:�^�:{D8�X�(�{�ߚg�|�m�8��U"T��g�,�Ƿ�/��,V-�Iw�"Z�o�kY#''__Q��J9�/�?��k�ރ�o_�-1��q��~a×��ʢ��rP�)�VDDĹ4�gM���V_�޽O�5�l��)�%��␀#�/�a��*P߰?��C���ܗ�.3hm�����Q1`A�X�4�:[��S�lll��yN*{�����/�
?*ݤ�/s�f_߉Fmޡi6BS��l�<�!��cw�n�~����\�G�j{�Ve�T�����v�ϭ����s,���Ļ��Gn�徎A�v��U�W	��$��ڞ�����sݾ��Ǫ*���&�F����x&0�!�]�P��5z����ۖvW���VZ�Z����� c�}��1W;���/���=�'=�!�ӱ��X8��m)-.���&��	�ը�hG���πv�źz����4���Q���u��q�.��C^jM��)g�r���ڶ�y�M
_�NN����604Ɋ��0�mT��Nl|�<�Z�|���7`ɫ1z���e� :��- [~���5��	�rB>N$�<�Y/��;���\ss�=w�����,g��e@��l˞()L0�)2�s��sP\���O�#�b��8�aڈ��L��G$Ҿ�&�j�d�}�0K�4���k4����ޱ���..�P��U��ۃV_v������mM�<�-�<�B�Dj���s�'�`��|��3��s��x�.5�ܙ��V�~���O7�n�����n��/�\���IEe��II	]��l�Rx)������:��NH�fܦ����O 	@��s�ޥ�78��ٟMN[����R6�9��MqyBy�����n��=%��]nͿ�6��]���ѬM�� ��U�����B+:(��##	s/�����XP(�_NBJQ���:�\����~��he>��=^��n���-#��}�=�\4���D���O������(=]6"b�!�1�� ��𿇦�y�r�>h]ë��j�_@`����2�F�ŗ�G8��S���&enz�*�9���MN��DC�/��m��x���'��?� �����ϣ�o���<H��Cb�Wm2%�e2�{�1��c�?��qmm�ot�"������{�
����"�N�d{�1Tp��Rg(�(��?��0Ke�K�����{@��&����NՖ�*JVs˒��t*�Ǔ'��2`yo�����b�cď��;U�ܴ��y���9����9� ���J�ɷ���p�KXUO�Ad{���:pܷ�
��WK�A��T�+�GE��Gq ]�����c�����G���<�g���vt��e�E�k!���s�iׇ��� f�����u���o`l_�� �y�R7�ө�� ��haN1��چ�~�j)ܯɑt�%����YYYװvbIB�m�����<=E��b���c)�rqe�w$���vFۼ���Ů��$/S~2@���s̯�Zϸ$Ґ�z���YS�� ;�h�H�8hTa]� {E7��T3��C�S�`;{�㉟���V���E���ԗ�0$�@�'Kr'k��|��l��h!+~]��'��*t��/T���>
t����%�ZJ�?"�L�nB��������h<����A��]�t�`���D��Z[��YX�Em1[z����넸B?������ݬ�9����<�;�.:�'�|<�EM�mE%ZstĚK������o^%�л�Zhܩ	��W<<�>�B�����/�I���5pᎭ���+�ާ���:�+F�y[��'⇁%���VS��|JMr�WX1��q��u ҋ���7o>�cjwi���4�wuY�38x~�|�k	�7}u�A0˲r>�fb��Q��`$���(ً�� �٩�p��<��~�(�:66��~�̿o`==��^�W9;�;�$�B�k6~zm^��˓]��m�����⍴�����@���tGB;M�?�Ɩ@!rx�)p��SzT����#o������9�" ��`_Q���F�!K�♖��3���z��-(���{�D&Ê�6����T	��oi���U�w�B��eq�{;n��!&3�
��Q��΂�w�|��о����/^(����W�z"�����j�o4{�}^���4o��g���Y}Y�V��c����c�
q��w;;��av^�}�D�����N_��豮�v�DTn�����U��m��(~
ss����{@����p�u�SKK|�Ws(�
u	g��ã�f���j�x<J�=�yd,�1##� �#.Ȫ�87�X~~~x�vbb"'���U�Av��:���=��z��ztMS4r�ʑ�L�v������O��_dV� z��Su�C����M}����}���p�/�22�P���߽{�>�x߽i�Ǐ��]�\a�{%iE;;;�N��;���=��M�|)J��z_��@���st^�YA#�Q~ݯ׼��wJO�td�-6Y�]������x�"���)c.����Dz��{W�g��Z>���xF$�aYkx����ɉ�~�PT���lF�p�G��ȁqd�Q�e������A�#�yGF�j6,I�����Xp������<>j��~0|{9W�j&č;_�=ؒ��k��Γ&��2@�OvՂ8�"�4�yw�}So?�'4�����z����a��Z�5�޻)Z��?�$�E+�g���Sjvs��A�cu_x��%Oy�������c�Eh]9У����]��;���ݚSQ�U�2�;n�3.����KH&{���Rѵz%\�,<x�!�z��Z��񩎾����u� ��WM�k�^ǘ�qȂΟW��8ha:Z::"[��k2Y��DQ����gNu_ٞ^�1>^�{�O3���cI��Wa:�~v[���ӧ�h���E��޷�O4�&������?V�dNl�-/?�����h	t�Q^>n�v��T�����Mj���ˆ��ox%�]N�mi�Rw��!ҡP<w���h������Ē�e����DK]ߢj����ӯw���n�����o/�s��ӎ�'��U�7�q�Goj��D��W�Hdj���k�?�D
YY�4V�Q\������O����[����):Z�5���<���&	����i�S�0ӻ4xk����I�M_ߘ��
+E<��g?�]di�Iב.�y�bܶ�dd����;e��;Q��c��M?����p���7o�h�NE���Nlߝ.LZ
`c�[��������F���m�m�츅X��2:V���&_�r��K7f���7r�\��(�|k�x.\UyK����˗����9䵭i��_2�ݻ�+���)n$'�,��hY�=��l9O,��5։H6��7a�F!!u�+���Tr���6�70ǆ����d�MQ �������nl�����oJz����=��_/�[[X����/s�����^����1JC�;N6D� ��J�`R��UWm��tї����M���d60O�Y��������㢑�.��8�>'�>�h���>T�3yO.<���
�}�89G[���n����P���M��1����K@�oW��Ҿg^�>EnPo����U�|b�C	^T6d�Āj������!k�/�Q�������$]�FZn���8���b��!�}}č�e�Eպ7E\��VΏ/�K�L��}�K�w��0b��l9�k��~U���rib,<9ِ�j'J�9beh�ҕ�T9!;ކĺDG�Z�Ba���2����yxx ��dd�f�ݹ�����k'd
4��P��<;]Վ"��$�g���:�g�+���öhDƴ�p�Y���b5��H��	.I���0��M���J�n�F��Z3��3M���׹�	B���&�8tX�?߁@���5r�n8b����P��v�2^HH�E��ЬP�Bi)�7�W=�;;;��Y)��Ѽ�0�xcl���ԧ�p�Y8��k��iʖ����ގ	�ro$���E���XXX�zHo���}��	pdbrq�M�+4T�)[�з�.`� �IdT����)��W1��Z86��5�
�����'f<���]B���������tb��[��*]�����I?~,,+�?����x�ݽ_�>wq��EI-�.`w9��e���;�uO�ߠ�(n[�E���r�ǋ��'�����o���=���l柕��]k8뇋���Pl�"#�!����̺m������Ĥ��w�����ý�A�[�=�m>�W]R�޶�"�.�?�����޺̹��^5X��x!V�N��Ӎ0����K���x`�v���o[\dF�x�#�;�jM�����e����jɇn���Baa{/)�b�`�:ƭ�J���o�� DJ��P������˖3�{�9C���L�BC���?}�[��廹��:[�{��΋%�Ț��M	>@e�K�T3�p0�c��}ً�G!W���ص��U��̗����<_����$mĈRٳs�o�KM��bXv!��.L*���оF�5�GXV�m9�y��������A�=n���l�B��]�����iy<�,,,��R�?6����U���zF�`���� ܫ1���f�7�e>��E��olD��T�F�RT|� �]�޳�C[�̽/�{���4�Wcq�m��;8&p
��>`��7�c�Zɫ�?%�3rPπ�c`�����Ir{χ�����ɫ����4q�Po���3����&����v������L����T��͏�Z��<�g��rmM�n��h�� ���W�CT|�V���c�VH h�Ɨ��Kӡ��.�t 	������5�Ff��fo,%cĺ�{�q�
�ߢ棻�mn�7U�?i���od?�� ù�$]�=?ݻPO���=�9�{7�D|,�:Z�#Z��ǉFʊ��]]�P�]Õ~$mZ�	��1n�V
X��K��v�E��U�4�wWF"g���~E�0�fe,z���������s�ԦvY廅��T�Gt��s��a�n��,l��il�� lbbb��]���'�����f�:Sw�⵻��k�Z���K��g����������3J���j'��8�����m��9B�@S����5�~�r�W:�)�RRR҇�zn)괫2rm�frr�}iT�<�_\RC`�ؔ�x�珻���\�aVgZ�ٹQ&!$�)��a�3�T+�i�E���Ϯ@�?XcB\%�p���=�}����i�����8�>��pm��>��y����3SıN�Mz�M7�8���bBl�����bAj?���|���{��t��ӧ��P���xHן��D�K�Pퟶ� ��@C�ާz|Bn�c&Nʮ�˸nO�ӗ�&I�Z3g�À �\}F�I�I���3RF�ޥ�x�E��3h933�u��q�%8�F�ɓ�]�)^����p�l���;��ʱ��ߤ�mzh��keꕬR�!w�J�x�#c��ϗu�?MO�O��aCy�f��a�">-,��4����卵�5�A_��P�R���5��R/��Rw{W��1��4�u	��ѿɸ�p�kD�2�0�2�_ej��䦾��"b���ח8WT�;Cy�L�ѻV#$Sr[��CK5��=�V�Y�eU��ʲl�?�h�n>�).GX�W_�U4{r������k7�쪆cȏ��ț��a!nTֱ|�����]&?_{��UPХ��~��(9�(�4���G�����|��h	�Q�������\\^PG۟/S �{ь�������wv�"M��28H���A���1{��w�!�J�k)�����[6���jf�z�B�.��\��c�Gr��ٷ���Q������ٙ��34��[��2_!�v��m}5�Q�?�?V$AFSRR�&1$+�v�Z�}�(-�EH��{��M�MP
Z��t-,(.�e�0'ot�tu�p˹{B���ݻ�Q�Pm`:""��޼�=ewU�<�*�<�ڰMNa�˸���4:2<�@��i���[-�͙�ڟ�}���$�M�Ԗ�ss�W���[�	
������Mue���s�>���c	X2?o}���@�i|`�t�=[�uv� �R�ҺF���^h��p`�7�HӪq#��r����Dc�QH�A�P_��V@�Jq#�к&�������G��);�����4:�HI�(�?*��jy��S����}�{YL>H~��i��qr�ϯ{�FR|�����hX%Ԏ���ߪ��n������8&mmm�������}}Ʈ�I�Ҽh�.�����o�`����zG�6���˗��&�F]1�v���#�W�-����ˮ�MG�c�$&O�mv�H�߫��S�����OSDzo�]�@F�'Ĥ�*ṂC�۝���Lfg�% �bW���dj�dg_���=�U�܎��Ғ�($ez?[ndBIBTt]d��6�cm-^z�Ń@i�p����Q==��w�&��TE\4�b�>wU~�ĥ>�޶�/�,����)�CF���jx'�� ����-�����і)4�_>���˰Ѳgw1*�S��J���R���N[�|����"�Cc��|Ϯ�F'[��\MB���������R��ɚ���ݗ�_��H.�=k�Z�-1��������O��b���%�%L�]��ƷKNBi�T\�S=�k�W����Y�b����r�����|%�0�UhqΔ�<�9X7���=�� �����N��v��ԙ�%k'��#+�)	@�L�ܔ�14�2��Hr��?�dߗ�GN�y�����r/�Z�J靃��k��r����%�MED�
f�7]����%���+���rG7Vi�<w(.ㇴ9��ˆH�X:;�#�{��X������#�� /A�u-��yl� ����H`A�y<�v)���v���c���1nP~���M^j͓�o���4���='g�Bur���4��4�^p������D�Gj �̒T��2}!�� "�a:����O*��/_�,����KP���Sz�'��"J�_jkmmmY�sW������7I�p&�l�$H�wU����\��ʛ�R����WGZV�-yÑ�	�O9�Y��EO5��`�8�j��KH�3;���*\�Q��ܶ�q���!`��ȩ"/�T���8�cSS���� #�.a�d�n�,/��oceZ]���F�4/��n���������O�5(:$Sv���a}��nA�B�C�a�I{^j�� �r��	������I���N�I�9��������o&8f�~������9u���U8�P��X4��D�[�6.?�J�����Y�t��2i�@��`����&ȩ�����5\�w�� S����;5T�VBqp����"C����M(;87T�#�T廉�&l�����g��R�l�gTWW�X&@MtN](�������
��T�߇���t� #9����{�7�l�a���#�B��]£����Q~������!PH��Y����k��'�=|��JI�i�y>��p��죽h(�`e���Mj��E�/0�%|��t=?���`T�U$�vb4]a:, j�~
%��4��t��#�圾��+�AR �-�S�mf�$&&�ſ!�G����Q)����]:%�VxY�Q�1�9�C�v�H�	���=���lKs��O߿ʇȉuF�߃��}��&�yi�H��@�#�%�b�+��פ�IdHSRR�M��W�Ww����W�������$�c������{|���2(R[;�U��J M�_�5L����	
Ȃ��k���Ϟ��>_�4��-(��7
�9�-����ʿ�<��M���rv�ͽ�I�
��^���`¹���n*}
,E8���)������8N�F:V�˸2
��l	���k�S5��������	�C���y��v�y��԰�GH���ɀ�ɨ�����}�^Ia"�3C��#u0��s�*b;��08����	�zW3/�=����R�ڭ���B�F��0��{�Y�|������-�`��$�*,���d�LJY��͐�����>��*K�1�74��K�|ގ���S)РE���)���z�",�~Q;��x��
bE܆��1ׇs�������˴V4b�w'�'R�(�C߬�s{��I��B�w�O�$'���W/�r���5w��y�h�k�%�f�{.���Gч!g\�C��c��M��F@�_��]e^ff��������|-B������������JH[&��u~ǍSL,�Ap�U g�vnq�@#����+��Ӗ���П������uU�cD���?\;Q G�\a�W�[��ߗ9���O��	h.v���۾�/CXE�?��B�,���T$���~تF�6��Gԝ,��4h�X��kY����D�h�M��=��\�΂�������њ4�P����	E����&��죆�u�h�n���Y����V�8a���z%� KG,y���6�����q=/?������������\Q<Pݞ��B0����I>:����#��fT�����Y'$\KE1֧��Fh��G�5P��OnUy�ڤ%-�9��Ɋ��4�=!����DO+#�0��j�a��	,�]�)�O�D�J�~t�-���`�����M�	�z���u���W�W���F �=b����D�$b���d��(?K[�0�i�nΰU;Om+�:�����RO������y�/Bc&RqL��T��^�8�iwi.�����+$�[;� 8��Ξ{n�h��m!mo޾�k��q+fko��J�Q���<;V�h	j�E���1/O�C9�q '��=ʻ=.ٸn&�������>X��r@U��+�|�9���1�vuw��4T6�͛7����JP	
�Rz����$����}����=���hR2�R����?9.��|��X�l��l��r�TI���Lb�������~���1[~ �@g���Ҫ��3�?�������)'�z�G�*ǋW��D�� @��%*���C�����^���w�����.���|ƙBA{hik�s�)~[s��3n�c���H�&�;�i�
����x�)J��p���/E	ra�}���
4(�Z��]��N�����d�r���yi�,�9��?y ���W2W�/��hDM	H�;�'��	�4
R��JQ4�ƝLH�{
(���D
�,��,칱��U���H�ﶼ�FG���ᕙ�_���yA�Z���n2��Jv?���F�z��˓�� 5��E��+t�A邛(%\��˙�i�`�L<��������A&M�h��B��z{{�hp+ّ������1��㲫��VA$�e��oC�ȈH()�?����^�	`�=�i��w5K��Raݎ������Q+��2�G��%)^6H�� ���2-\⎎�}\���#����M���z�l��ѫh�
�?U�D��+8؈�w��d�Q|� �s��"	�68ynKmz�N�4J�;[qY�]e�.Sn�aY�x�`D��*����MҶ��H��mg.�:N��B�ļ«e�O���>R�e1���:�0���O���)���
���5����Y�L�в������;���H7/�;4�Z��A#��d���)�e�8�[�����$��A)��5�3d�pps�bJ�P(�n����|��򧭃�$�Cn3���TY)(�����"�w?��{إ3�o�7Av��h]�M�������rb^2y?n�G:)ٜ�&��j
HP��}_�� |NG���X��Fm�ڧ��M��M�`ԃ���";U�K���ʪӧw#l]AOOo�hgJ�ځ4�����L_�>1ؔ��]���;;\�D�X��ؓ[�v�h�$����.�1��<s4�Hj���>:��3����Zp��t�2n >64Q9�j�ϵ껇E��\���@� Pf�A*�} kxm�mH��m)��$|]]U�>�N�\	ݦo�Ő�'�~K�-$ `�fͩ�>�RQ�g��g9��w�g�`f
���U@����D�Q+++�M���%�Q�ժ�h�h�p$����[� �n�����G<=F.0WGO�^��ۓL�u�߹P����i�l?�#�=���	��{��>��Jk8����M�D�x���}�up�1x��Y�xA�s�$s�f���x��&�W,������E�>��>V���[��h@��ᡐG}$��kE��}w�>3�Rࡑ�M�t`��eL�$�!�&L����wZ���7���L��d�7J2��7b����N�+������T��2�*(���e_B;�9��Y�H?㜦@�𚛛G��H�J�����CiR�3K겝�ү����fgAZ��ZO�I
�OK���[P6�&(A�b]C���yu_غF��tL}�ҟ`�2l����W������`��rGQ߇aB#������֍:!j��w�beܑO2�3>iQ����7�4%Ѻ��M8�︝�W_0�2ɜX�G%{�F/�a�ـ]� 8�Q�����ӓ>�2����kA��}����6ͥwf�J�f�����^�\�>`�����+z߬nD"d�>��N���Q
��.�z�ѵN����a�ԙ��[�A�X��Vx�N�d>(q�j>��+�س �JQ�4d�J�"M�~�����~|��8���}��Kc���A@M�n�ؾ|y�?���Y��~R�)�<�R��s�9�ƻ	��Z�I;h���Jϔ��&^�(U�L��O|��&�ϯ��/�ۋ۾�
>$t�ӧ4��E�­b���Z-�y��
����M�+�8pS2S�����V�����6�� �
�	q�B'����3�cX%@��F���u���F�ZS��JƔ]��F��l?§�r���H����Y^���O��cN�sg�"l�uh��]m۬��"C��8PAq1�e"����6�M�>�J0V��o�S��''��d=I��n����@��#䝪��G�pto�n��wr��l�>���F�(줞K)����e�g$�����^$ڟ)��x�9;��K/��	9%}��Bޤ��SpLN����2�\y���gf��>}z���+����ן/Pj��( \-�/���Q�5.��8�\�vw�^pJ��#�q����7ӚO�B�s�v٘���PK°���}��_���<B,���F&�C�����Lp�Y�Lv��ڋۿ�" �"�禧���@o�R�22�|"��9`���$o|HpK*�$M�v��X����$OrdK�E������\r�
DZ2�Y�88;������ ��S�+Wl�:�?�]8_��7�����C!]�ZWG�?<~��?,ɝljFw�M�����5\���z]{u�M��f�53���t����;�����Ecc�S��r�S��ɿT����w>�x=�YU~Vn{P��>�K�	5Mާ�AR��!�c�������_�g�ǝ�H��F�h�Bn$q a�W(@wr$yAZbϽA�7iiZ�,�d��į�]���������,��k��O��ߜ��w�'��d��\oA�����R�y�2��;�$�����Wf�K]]����c�#��0�p���<N\Nd����ϟ����5�.�����4%
;1)	��w(#�i=c����l���d�A�9�b7YXY�)��x�01��!��]���4��4(�#OՔ?b�?]��\q�E�#�PJq�L;� Fy��(Gh(��p�ϴ�x��H	q��[�O�7W�*����#��C	��ݣ�¤Q�G!d�U=D�eX�Fqy�`lPSQ�����r9ƾ��9J�ƀ�xǤ���n1i���	-����;s�W�:�G���9	R���^�s(��a�k�7t%k�~�Է�X��(�t�J������r�����)i,�gc.��W�9N�dwr{R;�>>�u�))�@<]�F�O����*���8OqIɝRО���n���冢 d�Ǧ��䔐�pP*Аb�������N���@�����}�%��kkkg��NGm�窭o+KK��RT|�]PP�q�LW�?E&Se@��2N�9@!�Meʭ8@4��q��z�e�����ى�}�v��>gB4$��+-����/��j=����������f��v�}qĚ/M�E�������<o�e+^j�͗r�ϟ=N��������?�
�������M� G�U�&��
�
9��Mj��>���}-s	�uM[\��XE旁�����n(�V�)��N�W(�ފ���f�9͉̈́���'�|:�t,/ =p�	Ў?Þ�:+ū^�q�h3��>2�J��VW���X{{�l�B6��CЮ�7��]EjmpA��Ii&��s��bTgڟ�Ƽ��������?�����.�>\J�}x.!��I�۷���i�>G�6����x-Sz�>�H]߉��ݥ~.���KCa��� &&1M[�z%��9��=�bbu�C9���o0�>��$r��75!_�l�u�I2,����rN�������.�6{^$�*3�������[Ʉ���j7��\\�q����͍`yLg��T���~�%RR՛���L�wA{��z���ϱKuw��MF��%���n�t�(�Ң�5�0~�B�� ��	���PWg��Y�U���@�s0&�܀@���"Op�"�c���U�����v��:���&��� �`H/��^�����h1��'n�@>u�?#EG85�g��	ص��|�'�g�s�gh�(�p���f��� �L�%���t,7uS�\���]�%qPB��ٳ������h�&U����,G2�
=��=/5�_�o�l~��P��@�]mO�#�>��������Dj��[#� 1�i��m'''-������D9��N���7
�$�K��׼�����$	���ԟ��Vj��
�j� R�n�UvP_}=B&�1[�S��8h���SO�z<D��G�~��HIK�* ��=J�L�0�$�Aٝ�YR`�G
�Ke�70�����#�8*8<���}���* �4� �����a�=�_3�]�9`>ǭq�h�K�舺��K�u���{�$y \���A�w�Lq��9
���_z�&*�J���4bf8C�`��F�[H�S�-(I�D�hn��P��(=B���{�<mW�����_���=��WT\iۙv�MTeK��P�7yȫ��Kם3h4�o�o'�kN����T,���.��Cϋ���Mn;�r�p�o F!q\||#�e��Em�\��ޥ�C�F����,9��>��S_sJb�?U�۴����)ߐ�j�5��W'ud�(I%�[��gg�H�����ZM�>Ai����W�m�͟�n����>�o�M��]�~�����/�s��'p��/��'����-D��ƃ���+PZQQQ�)�쾐Z�8�ׯ_τ2F�~z��>����r�eA�:X<�YK���6���3x���{u�:����-j��7�� ����bo��jh�b*B\Z̘�j-9Xr*z����hG�ׅR�&>=o|�I�t�	\W�U'���+W*�4�������23/���y:)JK;�kh2ƈr[;m:���~�3W|o,ba<`k䟆��������*J6 $)��Dv?ò�O������W�4焆���Qr臮�Z�׈��*��2�����p�1\,����Po����<A�؟��載̷�G^�>�T&yV�U9�Kك��Xx�aPƴt�����:�H��	�÷�O�WW���y�xߞ��������^!""j��L766֏1Z;!!!<{1��-_���apd��'+��[v�)ǜCŬll���t�
[���@�K����*�eQ
�>=�����n.���.��k�Q�222;�Aj��?�����\Q�W�x�~�aĺ}��9[Y�	�~S\��5��e��xxvֈy���������k�`��;�$ZE|�F*�_zz�¯��t��o�|
��!%'�'7j��͚���0kӆ#з������x�| WMMt��ә*Գ���[[!ZE2ZZZH9�hU<�������`s���Zm�%��npp�����n��Ga����
/�*�4v���g~����M�i��RaA��fE�Z���������䁟?%r7����u3
Q���!%�eIU�Z���k�U܀r�*:�(��hw.AA*ȁ,Z8ծ3��`�[ P��b��Nh��f�8DMj*wpr��j��E�j`̖�uRRvc��Н��ү饞�C�eN�8����8��tY[H��i�3�/4� U9��"e��؂�����CE(x����B���u���"���m�V"�?����#��������lF�L��!|a�=^#N*N��w�]��w���LV]�a���p��q-�f��x���d-Wt�Prς��Ǐ�2�पOv�K��
�ݽ;Ow9��|D6������ZQxcʸ⹥e��tX萯B����2S4��E	k��������=�������8h����Ϗ^x�f�T������dd��+�RR"�|��>H��𾬬�`j�1	��g����;��y���k������p}�䝋xv����-w�2�0e��w|�%��LL,��ijn�!��B���� �(�S&�CE�H��Mȼl�64�k
���vh6)��G�y�c���!�����+B������]Vde�B�=CVB��P��(�d����u���^������s�뾮�����>�?TR��\�ؚ���u{{^�z��<x��Iϟ�޽̛I�2�R��x�]c���y�vr��T�I7�Oʇ|���Tml8���&&ʼ���� 5ԑ�����%4s=��WRr�b�N��/�Q��80��-�Y&�~)��������k(�� ���1�����%��[���"Y�r�z{U=z���7D�]�u�-�mε�2�j���2�|R9�nݺe���&)+����Δ��\�@9����ۛ�Ƒ�����,P����s��>~�|R�#Ny�I�ʭ[T���XAM��Ƽ������@R�IR""f?[�d�a����J�i�u<#�{�n�E�d�"[�N���{��ҷ�#�І�pT��=�[�
:�JM�$�A �# �/�Bxa�U�G�n�`aa����	��Wf݇�%<�X.++����9*�磤���fK�}���y�*J
�flM�k�R�V������A���<
�
�!�K��L5�|:� �����yysّ>�0���R4��4.3�r�!Tk˛#�)D�o�훜$��!�4,��YTT4ͼ�FgC�tt���թ*
qc��>�V�u��!��׶�*��'Zx�#y>�~!���NN����ѐ���10��=2��̠����|��V���wj�^����vlZ}i����8	OZ-��\%���WH����E���Ϯ�����R�i*�Br�}JO�l���B��
?
�x��������1/��cN=��1U���vU��T�VuMM;D��P|����ׯ��Bxg4���CUy��jI��	�o����Z�w��)���҇�!��a�\�w�Ut�U�����RSS�	�Έ��*Trs������zKX?A\8���j����$ۋ��j��|(�Ш(|��$q(SSSQii��,���rJ����-�,&�`T�%�C9���U:C�O1hK��w�șȹ�������<V�J����%C��S�����������u�AI%$�C�������(��CM�\��"tx�4��7q_?�Z&��=[���RBh�ǥ:�	xP�<��
����Xjǈ�۰�;)�#l/�jX>����Q�ƥ�ka� ����566&R����OF~�!���[�c���od��l�^�����M^���TY�->��� �j�%R���z&&&����ꆚ:)��d:�K���V�;�WIq[���n2�8�����/�T�y��XE@[�∁�0G�п� ��q��}��Qqss��;o^AC~`�aN�`�ޞ��}���H/TҸ,3	P��|�����P(}�?�O&�-�^�ꨮ_>mE�����p�1n������;�x;!ee��wH���c�oH��45�'J1����ݪ#ի&`�}������\6JJJ-�����yqO5l�q��M��l1�B������0
1���5O�~��"3�.����.A�!P���r�/�/_f�!`қq�6���M�p�����3�
J��rCC1ќ�v�(��d
&o�MՏ�?�@���&����u���+��9���W^E����̗/_��A�~5��&^����[�в�����P:�[�SO��f�>>�[
� ���Ah�Y��/M��<^\Z
y�N�Đ?x��&��Ǐ��:7�(b3�?�ܼy30=��}��HEUu��{�����������(����j�����y*�����ѹVu�РD���
�VӃ����\WP�x�G���ߏq� -�g�A�L\�"�)�PX����TZZ
@�����JZ������m{5~������Y�\���8�3O\ƙcnݻ�]j� �&B3T/,����	}'���Ԁ��?2r�b���������H��93HƧG���� i�|�I�!����/�q����KKc���j���Q?�
V�5�j��H�V�S B|�b��� ��|�S8n$y�@���K���塞@�`��u���QG�?w�--��K�7Wi����"������UUC����=MI	���E���%����e?��E��{zsj���5�+�&R�w.��<�����Ͽ;��' �.-���4�VP���ͦz�J.���Rrv�8���Y���w���DAIAwrf��C��g�k~>*ʎ�����"��odDrɽ�/uFMm�E�4>>�+�Sԗ�5�Z�G�t;{�H��r{�<�vMj>>�:�~�-Bb�V�-�kT�� �g���q\�,��-�Qa����D
�\��ދ���v/�����I�\'#t@�K
��U���"�GW���9�م���G��?�TA�F#c�.3�^]]u�-7(�� ���8������=�6�e�����h�v�����\��A���	g���k��Z���u޷ �>I�������}����d�L�y��+���D�b�����Aω(p�^a{�����,���`�2B"�;vv���-�ܯU�I��%��p���N��?.�"6��l�&��H�Rl???ZF�8.9��B��.`�Y��(�A������ڿyC�����Sc�H�Y����͖�W��t��,ԓ��M!��>	(+��j��zF^@͊���������;��}����"�����JI;;>~��(h�����k��t���h-3s��H�Vż(�����.K�;�f.�|����<?�����W�L�jW�4���߶��SW�b�9��&Jg3�l�WLL�/p�2{*�P1,�`r!��?�)�s���]����û����w����	$�L��`p� �M� ��|��H����X�d¶�uc�mc?<�{�E��2T��H�� �Ʒoh8	@4���D�!�V�rY$�)�#�>�y���<?[�x�<˓CGx����,-P�UOP$��z��~0�Т�JR�Ka�)|��[�q���G�3�$r%{{ZwXO��s�
&Xy6���- �s d��h�#����	���9�\ _ ���>�$�y��wCT%���h�?��~vYLY� F�%�t���?���?j˺�%ϊ%�I�q3"�z#�g�<v�k�>2��P��F�<M�(�0�ckq<����,i�+�>B6����P���,�{籱��G��\/�x̡#1��w�.k�R²]���=�2�i��/�ݻH|\���:vh����%���p��A��N�o;��|�9�g`gs���-�r�����"ސ��Q�/��~�d�B�����B������y�0���ZSc\�}M(� 2 =	���h./�3��+BKط��p��i%�N�0ؼ�� E���O��e[':���\p�j}�]��|
�ې����)	J՟���6��f��2��	�]��	I�	#o��fPb�-́ybPBt�RO|�w1X>�A�Yi������~GV�&'{��b@��piB̅�KHغ�V}x��
���k��P�{3���LbUΕ4��h�Ԙ��	Ǫ$G6��W��;��Dr�ǉA̚@��t��'�<�����w�I��3��""803d��t�32�kE���d�IqCT������qMʘ���>�%�6�⯆�_{L{4Evh����}�V0d8(�6I�_[�L��ӡ���e��pe5}�(/4^Aơ�8��lml�V��BHg8��0��(��i�(À�%R&pĪ/+E>�yDk~�ȿs�72�����d��c��{��[�K��MMd���1���m��jhH_��S	I�U9�߽s�:f�>�N�3���Vs++MU\	f�P�_�OH����윜lhQ���<�s	�I������u��h��ZpEW����5������=L�diU9�a���iL$>RFZų/& ��_R�y*)6��b����<���)��1333�T��IO��Pi��*z���NτT����\� �b�/"�4��9� ������.���w#�}@�NF�J����]\�K�)8q��u�9��֘ -��L�r����!��\�62w5����$P\p������[�ڑ�(��c� 8U.ދl=���5�U ��$���j����A~]�y2K���z��ctG�|�W^.ĵ�Ƌa_DKm�����h&ޚ���)@�^mm���9��xx8��1�Y��e)��q��x\�h
P*��TT9EE<�3�y4M!e`���^�X��X���ӗ��~��5�3�pN9V�t-�o�bw�㼤��fv����:�6?�[�A����6&3��%v�[M��ZC����sww(�L�e�V�9�鏫��X(�B
У�;�B��e�N�R?Ev���� )��ө��V��-	�����%�ٷb$X�d�����"
�7!�Fo,�^��� o����۲���a1N<�O��X������NvI	�����N�=��Ks�����H�]
��y��T�o�,˒g�������y���qkos��J���v�0���SNNNv�����8M��6����F�=@Ů�D;-�
���[?�<��`J�Z���]�yg�'���L���K���2�� ���/Y���8��R��í� ��5qLB���a����<�2d$m�����W�L�}
mV���ߪ�w'��B<hc���V��ި5r���`f��>=(�q��i�s���t�Y&]Eh��ܹJ8��I�J�&&&�圠�E�A~�w�Ҩ��<�������z/�w�Q$r(��zk������[�,�b=R�:Ypx ��x����4E�ng���# )1N:HSw��Ǭ�������A��{���ʘ��5?�7�7�M]f�H��"�1^7x��|��~�i
��!)L���
z�	/T�y:N6Н�4����~����uH�:#�~ղg���� 6w��������e���p���=�	��	��5&[���*���6�X6\u�)v(�ӻ�\]�>��ͪ\Z����	8S&>�]�CH�ݯ�fT200�+J�rY+���1+*�:\��{nh~G'��H����F�$��@�"~�����1��4I��V�a�{�v�����76T��$�Hm�)��h@M�_t��Ԃ�#N�,���� 3IW"8��hh�Gpv4e\&���3??_w0��~��Oh�kvN��ޚ��EjZڽ�p�B�G��R���..Vps�bm��D�2��Kc�廷��mbF�����~,���'Zh=H����da���C�����k^I�m��D��t�渲xJYcE'�Fn������+�4��*4���scO��!�Z�}���(�J���]�ɵ[��j]:���2^Ȓ����?���t%�Uv2G�7w��V����KH�(�|	�[B��h�E�]�h�Y�h�5z����q�D����g���C�3֝�Pl�6cb5&�������QT�o��c?R��~�{� eb�៫X2�D<d���'�,��1ui8Y�(����RB�`�&q����i��dM�v�zF��t��h�7K^���zQ^\�rץ���Ӎ��H���zz�I)�!둵��%4e�4��u�X?�r�?Y�4l���X=E(��]���O�&]�h>;u����^�`�%Bh�sq�������?��O��	isg��kɬ�SRRj\m�o�4�>���6�a��"��*���p#�����$�f�2�����N�S��d�0	�(��oL���e2���%�ߴj��H0T�Q~�X?��5���X�:�]ͽ������~���2�qr�� ���_��gh��f�2d� �\V�{�|��n���3����J��'���煽2�,+����pZ
Q�!�D���5?� }��"|��Xt��WOp�����U���B1z�4�ϬV�����og{C�7�\b>���Zq��b�Ca���J�~�6�r��u�^�"�����S3�q�[6��>��m�e��ݻ�*����Z	K�������6����/{�3��Tt�W4$��D!k��Ɋ�P��� Ey8�+ikk����Yq�exg��-��|ƦN�4�$�o�j'�{�5>M!�=�\�Y�p�bk	r��N��0��c��/(��q b�&3O�Z�TE���.�����d2.p-bx$%i$�]��ȟ�=���ܑ�p<<<����j�
�n[r?�/+�K�b~M �p��^o�|�߹���߼�b/5�Ύ�ݾp�h_��}�	����o���(�tRRfEH�F��AcNm��p뚏����-��h�^�k}<x�	8D�I�����i(�/o���=�^G�R�!��,JKX��yv���0���+�|��1�x���	����d���,ͱ�&����/���۵VX�D4��VLl����~�G�~=paE�g����uӥ�:�N�E�¯_�|�Gѥ��{_�c��6�f�����.Y�10�X���N�~�MQ �����/a��-ݒS1���/99�����F��)&?�%px|~{���=USS�gqɾ����o߾�ן�RF(��2?�@T*��#�E�f`��G����?���\��ƪ�ޮ���>Ƚ��	ﮌ�9J���p����f����l�e���pD2D�� �6��F;��0I���U����`jtIYY����k�n����W���qh�U��bEҺ��l>�,�mn����Y�Ym3-b���0gx�ڟ�߳90]o��;::�����BӴy>qj�B30t����~�q�6"����7ػ.g��_�������]E�k�$�Z�$��W�C7�VU�	!P�6* �c��Ç���=�F�v����v�Q4�}^�~�7�>�)5����G����K�ɞ�J*�8=��?��'k'�p�ݡ �=2��x$�r`>��G18���x�1Ra��ٳ��T&�&���oE �A�a��T����8�4?Eo��?_�^�!w���������KF�s-⭏?�E��-��S;���?�pZ5P��UZ\Q�����l���j��$G�V�[�1�Ai�m���ׯ_U�(N��c�]uf�v�����Mx[PO���6��o�>��O�j��������O�<6E�pb|$h	� �G%��9Փ����Cut��,�׭���<��Ťu�]q�\.�b��{�Ifv���s�g:t��=��	��>%^���&��6��,�&O�^�������\�y�9�
�ʈY0������cQ禿���∤6w�޼!mp�Vs��]P24��/�����>^�T�w�^�:�tKB �����'i,�O�|ϗ'a⃌I$�������f������z�F�{��q����{Y6'���#(<h�z�o��6�.�L���+M
�Vg;�Q����������k�ԂBe����������98���$>F�`�(l����I�	-��ᡮ�����ޢ�޳x�TתF���\[[��n�����RO��9�����\C�+�%p��Fw�JNJ-�2�4!I�������Z+����D��G;��nGk���\�WE?|7�q!��\I9�&j�d䕮k����0���]�4��xxy�T��.ކd�PJW(d���&��7=���g':)IZ���	�Y�A'�\A\A��4�i[nY��n���}��↳���Bv�z�F�F�pSW�����f���4�*��l���dl�}�"ͽ�\��������`֩�r����0;�����͒!>�ԝ��d�,������	���6��QM T��wS�~��Q���~M�q읓Y=�,I�I��\iF�ha9��A��[�bbbn`+fc�z"?$'S�y�R���@��S�:�(6�����ƃ����se���#B���7��qё\��}=�m?T<6n�y����.���R�-�f��	O�I�<Z�TF���pjL����Ĺ��Y>$V�B���N�3?C���ͪ��?�ehd䌗Z��ʦ+����&T:��D�Ê"�q�!}SS���֖�ʒ������ ݙ�á|���G�N	,���`�_v�ɒXR���� ��|6�l�.�-9�X��ѿ[�	��K���:q2x��N�K#\yRP8��������1���n������a;񩿐����qG�OW%P��p+e��n}f�G3�.-/�O��L�� �U0�4L�E����l�LM����P�x���̱į�S�R � -#�'����e͖��W���;�>�K��615ퟚ��L�E�b"FV���2cc/ӵ[�i,d��ʟ�INz�}�ul���ŗ��D�~�oH����8��2E��� ʭob�-w/����&x�/�����F;T4Rk-�o�$�t����@�u���&�jo�T��C�f͂��zۻІD��B$q��8�N	2��Y\i����VV�67]�0�Yr�VʋF�A3����r	v�����Po���'�����N666�o�(}gJNMMum�2���)�$� ��ܜ���V{K���4��^��)�R\��y���qW˲~b����8�=I�ng@���W����＝�c��';����vp��B(�,'D�[# ���*A��K�OB�8�L��5Z�I��#ږ����gq�b�������:_�m�����P��W��dd�2k�~���Zt�Y��ښm�Z�u���2���N��j��w�-�/Z��VB~3�g��	����M��SV��	�B�Ҝ�Ĳ���|	�rw��#��T1�Vsο�
Cv��-!�B��t���咊8'gÒ��a�v���[?4��P�t����ڀ`(�`��%�Ɯj�g��j}�VD80F�η��z�Ǆ��AV��>
����}}o4t�.���-6t���{�v��+(���	������Ň���N� }��!	�*N�1��u�E~y�Ɓ���ŔU�ެB�"EY֘l����DU\�t��iQ��Ph���w�i_ț	���c䶤�a����2\c�x�Å�ۊz��	B!-J$�B�H�*ώ�n����?��t)����^Q]� ,,l`�����_{qu����Q��_>��ʮ�N����~�7�Fҥ��j�,�JJ�1������d���r� s�M�j�?`j��'��7+[آ�Q��?�����kVV���#๯tl�up�k	Ė�(h�^SL5<�Ņ�����4��T�����F�o)�<S�kqc�3����������qr�v��$]:����+6��O}���ێQRj�@�3���ϥ:�M8�/�c�כ����I
'���I��SWS��.x���`�$ "''��Crxh�����.����u�xW�v��+�y:-�<�JR��&�M�[�]�v���cK=}ABBb�1�HKK�%�Y��� �;\f�D?���El,�<�PF�x���L���;Js�5�����H��?)*��i�%�|�������� (n���.�!F����ބJ���++�d��	I�ތ�C.��ޙ�������߽���	3UU4:�\��UO����p�8����I�{<�\��e9��~>�2��e1���Z:��E��Pq�q�*r�(?��hS���95I�}�������ݐ��3֘�S�O�B�{Q/a������M]oU����c�=���H|ٮ88؆Έ�^\��ۘ���#���O��~�
D�P��2�l$��/���+	X�o����J������ӡ������i�r���$�>#R���2�4�����w`O�z�z(�@z6��eݏg�Yf!��W}��gK�z�n��v:����P��DY�r�g<���6��Q���?,�j�d�o�����A�K-���bP]|X?A����A��g�uu�Ѵ�,�k2����E{J����a�~�Jy}��}��]Hצ�u�!��e��m���sr�v�~F\؄q��ݮ�%��Ƿ�2�J��r�&���z�����s�[*s�Ų�2;gg�z_��@�[FC3�������^�� ��KqNMMM�IϹ�Ď��+e�|�O��ⳎqW���=9i��3Dڥ���]t�0����E�r0��`
Pώ��L�3SR���^f}�ȊC-`ȝ�=u���~J�����b$zo�S����j�l�bW 6��A�t��nDr:%���#�R�o!�0	%�222�=S�<B���L���L1Nc~>���=�����sF#}}�Z�y�%%%��P
(�Ės$�٣�+g���Lצn2X�濚�[�(ꦟ�%F  �b�7�7�\�eȸ����i��c��(���o�:�
s�/�Bl�m��Nۚ���ݻ����W�����<{�{.6
/�c���J��I��7��/Ϋ��t���*W�\��v�*����_�'/Ǩ�A�ʞ�I�V=��b�͟�����#��w���qrbb�C�{��q�g�*��$ءS�v������D���Y��Y��&��h�o����{p�q�\M��
jԶ����ᗲғ�9���z�ǅ`���Ǔ��5k:���塒��z�Ⱥ��w/66�����m�S��	*��#fcg�;l���v�tH���aې�����{UF���f����k��T
�k<�SLȏ؃Fem$��)�[nԡ^^\��D���Ӌ�Oz��
F���C��bl���edh�\�2}�y�u��rCfw}�H�!�P�~����a4�	Uz��Zl�w���g>�$�t�)I��g�%�ߧ�y���I�Z�"�l�[R�_X���-4�[nCRBB����Neu��6;j��p���Դ4�����Ol�����{���w�(sV�![�Ѧ�, @tV�����S����~�:�x�6VJ� _cִ��(�O	���1�`|~�ؿ�`qD��'�a�@�x�{yMYI���>²V�!���,x�l��I����L���U�O����Lk�S��ˠA<���,��t2�
���G}���F�r�b�?���IYO�"]�^���:hhݽt����#n�
'GG3��g����y��^�O�o!�b�YjQ���9���~j��,OԖ����g��o�j5��A�i�r������@�Z~ˆb'������S�s��1v�?�1��m�C�0@�Ox���c�����4�.�f����#�<�LZ&G����Z2��')��r��-U#��.�;`��%��:���ed���t���䦒�����ʢ��D���VܹAd;]B��~�i�G�FkL�&D	�lہz�
tPƤ�|)��-�hkk[��������Nz%�����E*P\����ހӇ������x/)���\�-�ȑ���^9�wK\_���M�>���Ƣ!�s��
>BeY3�|U[�W�Q�������oVr`�!B�dL�Ŏ�u�<�����/�I����S��XbRŖ%���F&�J���F����{3k.Ѿ�4TTTOm�|�V��U+k���?���� *"B*��5N�Ug�).!������+�	�Ht���Vt���m�Z�A���_�p֐?��$wh&���s}[aD�G�|�j���w����[���QHD��@�V8�$X�s�M��			-_i��'��~���:��N�.~�K����_hƚ�SLmXD\R�>��mvK��' �C���2S�v���b/rs����B��Yτܛ씸fba!O�;�IpX<��Ӥ݉8������_̅����Q��
\�h4e���,�tk��$A�A��z�9�al=Wǽ�����j߇�`tH6���D�5#��@�K1�]Zg�'ȱ?�",.+��Q����^yy+?iM��Ņ�q���M�|fB��}�K���	&�"g�Q&i��Pʣ������.��Z���vww�1�<��%�5�clL�t8T�
Hrm��i��"��A��Ʀ��s��0Ɍ���"��� ��,�u�u�UhU�r�=���g�h�������}��[��!�6�K!��`}�+cbm�HQ�¦��ZHZ���OڿL^�pt]�C��ӣU��ͦ�dRF���V��I�#r��ȃz�����j�C����]EII�Z�`��D�J�����5�RM�^�~|Z�WX���Á�a{��6�C��B�9�)d�#B�~��,?�o�y�d���o�k��)l� +�azD������Fh˟P�	���_�0L�Y����%"":�R���M���X���!�oPz��h̩]����r렋ZK�p��=��9�|��+Qˁ����@c]K�dR	i�w,-Q 2`Wv��r)YC��TTU/���c|�������\��Ujs�~�S�W�VA�%�1�uI�驽�(b��G��K����B��]ɝ���	8�h�Tĝ�3�t�����h	��'z���b��u�}� 3���W0�d:��l����Gk]X�s��%@�Gܕ"�jnn�>fË蘿��1�P����J$��۷��Ґ#u��I��+�%������K�'Yg���A���ed�����x����V��D��_5�C�]]�8� ����n���`�˱��T��;�{x���GEx
����^;��R��	
�+����I���W+:5���
���Y�A�~c��a>�8CFiO�j�4f�d�/���^���h����6�Jd�Dy��� ��ތ�!{=����b���H���&�����:���IH*	�Q�wtt���Y<@n�,B��h�����<}`rd��oG��(!�J�����^�%TY���5�ǯ�����6Vŀ@�sOϩ��P��������Be0fz�!�S��ӗ���_>-|�/��f�.h�.&cr��L����Φ�t�������2������>�Lh]�E@�2^��#(�θ��?������i�͏�mPo<V�#p�_N�EE��&c�y#=r�7�ߍ�N���7���T��m�S**H�+$'gn��f�k9�������l�����'�(jĶ��IY�eQ�\/l]�n�츛��wE�O9V�<Aj���,Lj��r �p6L�:+��n�D�y_�H�������k���˽���鉚�<�����6�uPSR��@)�Z��L�#�+d��ϸ,a�^�w��V�=9u�2%��Ѡ�����p� �"�zvMT�������r!/�',���qdA��O|�j�o�t�ױ��5H�(6B̏�������JP����(1B*�8
^R�D�0\�jy��Y���ٺ�����r��L�k��T�
j�������W.���1ה?C�2����GSF���\V���x,|p_�x�جT+��O}�����3����`��F8���1�R��;�����w���-ʋ{"da����jdaG�8�m�d��Pgf2s-د"�***�߲(�s@A�O80!M�Z<�����y��T�5
�#�����x�pM�9�F��~�+����$���4�s͙}?b�7�Z!�~������*Z]� �gD��L��?��w��sc2l��(*�gC�А��<!�S�h�1�Z�X-+�V���������޾�#6����9J�XF��s;�½��%�\�gE�q�~�m�X�?��F�*����>�&�<��Êl�s�h�_��ŃM�����ܹs�U�H@.�Ԙ�oJ�xYWN+%�e��d/B+�=C8�*��MoW�����@�����%l,T������'9�j�͇Ŏ��M��	�"��b{z�Wgd�� Tx՟���h��Z�-��f.u����+����X�}��lqeEIE��H	����^=G���+�M���h�����t���h�����I�`~KF�>9���k���'w/���lS]]��֯q[5��{�*m��ý��W)v�e�T(ǎ7��W|���x�7��\�#�Ǘ�}W+#��z�	�څ_�+�{�#�#SS�w��w��E�~�Ix[���� �|���h;��g�m3P�{F��He\��ٙ�d�\g�����l�`��ן��o,/C��=n:4�@GZ#`�:T�T��l#����( ����"5�Ϸ6�1����MU�2�[�����t^��Q��З\G�x���ם������5M͹�׮|����/il��e�������GYYmjj:6ږ3Q����〺��~,�B qrr��R���2�l|�v�X�!��j�q뽶�N��t{��Fs�/C�;]�����(Q^?n^�g+nt�SűܫZ�DD�-�����ɖ��Fo������o��fͻ�*
���vU��&�_J3�y��(�������Oc��*�py��Yp�}Ĩ�y����CII�����m�Q�F�gW���%p,����tV���{p�Eٱ���:�ݏu�ۇ�)�?���!췤.��Z�mU�m�B�] gI�����_ ���圇���g�iD6*~�����Q�ϕ?0=G!�Tϟ?��8�lPfr�d(
Y�
�1l��p�NI.X��z�=�80
n�42�sO	P��5��]���_VZ��XC�R���3��?x�&��.ks�ܣ�4M٣���R	K�&e%_��D
ԖZ'��I�*'���fff��\U��<!�0P((d�mp�B��;G�ӽ��N�S��dSd�{��е\g#�{��o�����o�ϭb>T��v��B�H����J�E�DL���"�'4�����j�ff�U�	����VGg'�4�N��+A�ݜ��#;��֪j�ԋZ�ۭ���j�fgF,n��e� ��V�G�R�{���^jYj�����1�f.5>�{{��rz����&l��t_��I󖎎:����7��m&��ϱ/R`B>~�XTeʫ�˱؟�@ixmUom���ϔj/*+[:�-,,���	I[tp�Ґ:���LS�׷����y�+
$d�!���q�� =B��ҟF�R��2N�y�^��e��6�������;�NƇ1��_��z.��ɬ���a�ht0���.�!�h��v*=(L�[�����**�ʸ���r{3�F����+d-�pO��xv`����\�
�a������'X�{�DG��*�ٿ���DnV����|�=�&��6�HE��[.�d���m�[V���V�<��F	v��W�.��L�R6 �"Pm���7�r��+�+���n/��G�����W֊�̖���Wܼ�;��f�{�,O*Y�մM�<�V�/�\aS��3V�5�Z�����Շ.��W�>���}q�����>���X⭙�#ڐ��'C�C'����~%^==���z��]�g>��o�	����D��Efo�;qmt42<�Ns��.
��	��(:����(�|��O�<���k�Q��z���<V�^L��W��׎2_`5~��HC��̟	���T8��M\�,t��*�_H�o�������^��G\=��ꬩU''A����Yt�Fv�A4��Swjnݺu ���{_�\LSk�k d��]q�g�L�B��(udZf���<M<�z�W��[MIV�]ɂ�F��XEX<rw��V'�Sz��o�hH�(���8c���.=п�����I�7_z��bq�l�|��$2^�l2���x�ki�=ǧ�.	D?�zyz��>�}�"��ģ�6[�m�U�R>>5��Zk�4����:htH8�kzL�c��H�m���K��÷}8�< �t����F]�z�so�����`V��ɇY>�|�6
mY�%Q��hᦖNu�wo998,����8R����R��A��NY��W՚��JMf���*s�+u���N\��t8��CU����K�"X��_�'�_O����
:w��[C�����jj���6�q���>��ѣ������&Z��/����h}<��.S��_���<�.SM���+#W�5�(^i�|�!�epxu�7���tW8��
�ؽ}FlJ8T�F���	��P���_�c���ڇ�K�²޴�^5'�{��t���9�8W�6��˼W���*��Չ���,c:��Kz��~�+,XNw���\g��ҥ�vv܏��\�E��	'���������#���
Ov=�/b�������C��G�P/D�yy�6����f�s�_��9y�i��R*W����Ho4g�Qa�^J�}����#O.y���|�{b��>�a�|���H�W�F�c2,<<�7n��8C���~C�kk�$��Mk�?�Ǐ5��NiYY�NH`�.������q�y_q�:y�x����x�yck+?��q��3�n͜ʴ����$p�76�c:�v�u�a�I�&)))J�ҩ���x�����л���>_˿�z��ϼ����9.�VǺ�Y�Y�_f*�2L�rv�sE~�'c��3�7��溺VJ����<rD��T��e���8�^|��(�r�r�?Wy����l�4P�y����W��~�����kEm���+!�(��]�~��_	z���x_X!�:'��4�Mj������L��&��WW���ӊ*^ӎ
R�d^�F&��h��d��W-�Ȣ"�����v}�XȝH�}k 
������	���ym~��%�����Ӥ�xi�]8.3ˮ7���o�|�eF�6��~L5O�^��z�M�<o_������sӻ����E#��)k%��1���[N���h���V�'�r��eW?�{8/��j�^�����A̭�޲5����WKN�_5�&$44G!��4������<�o�E�8l�0u�f�pb�}��ʎ�f����<�1@�X�����/���PFf㩗pcv[�%�1�~�8�]n��o3����2N^)2�����(�E��ͳ�h��+E��`|����s�bfU�.�u5F�8}&�b~�R��vʽ4	��W��N?)��Ѯ�"��������j�"�E6�
t�)C+�k���əs����J������ U3	��cD���Y���Ƹ�zh����g�t�5/ru�,��ja��t�d�Oke,�m�������Ŕ���k�t(W^�"�O����ʚ�"P�=����D�Dw���ݻ��G��ĕ*�M�O0<55��'�ʕfv$��*FF/fߪ�M.u�u2�}����e�YS��7g*��Dhii�ʏ�{	�V�K�o
�Δ-������	���Ń�ߊ�=N(3�O�_ޚu��ܜ9|�־+������e���̅��1�'�.kVs�x�͗����$&6XΟ��8TB#�8:���YXJ��k�Q�l�E�ɭ����90<|||��A�pq��*O(c��-qΟ�K�_�0nU�r�rN]mhhhDttۛ;m�U6!�r�)��겑�Z=��@u�����+���m��t�ͯM^�,���pV�`#���k�"2�h��l�'��b���lzU�w������«K��^T�.|�\m~7ʚ�"!m�R�d��pHx��S���m����M��6 �c��8X


��W>���y<w"���rWQAZ��2���%G+�H�ް�C�P�9=\a��0�Y�Ɓ~�,lHhݿ�N��~�X���F�]���T�2y�ū�I�t(Ӱ�^?��g}+`�s&�u�ܢ����d?��<�|al��b="{�"�2y�T��&��^y�lϱ��#�O��{���unQczzzWy#�J�ӷF����VmL�,k]�Kjnb���'��
�X~!
�(��kQw��r�N�Ыa�u����S�OxVo�Ɲ�%1;J+��T;����]�����%��?����.P�+F������;4Hh�l�)_��S���UT�Q�/�"���t#�"�%���Rҍ !�t#�  (J��� ��-�%]��p��w�wg����c_|\0��'֚�+�Ss�TW5���q��T�n�Me\�����<&Ù�,�����4�M\Ӹ���|:�ﱬ����(J�����E^��BCCܸ�axu*���ɒ��9�!��@�����_�X�i�����\޾�̟�~��q`W��Y����C�1| �f�4#��l��vڙ�
�~���QM�467�Etb�Tڢ���gW#�֮v��a���^�%a�o�F��X]���Ctllr�����EUNp��1M-���B\��Ow�mQ�e�c��d�}�6u�5K��TSB��2�����|e0�Y]��;��3�h�`��%��'#3�݀[.Bђ��D/�I�1��lB*Du�h;#���K=��uF�V~��!~��1
�"���;B���Cu�O��}㚪1'�z���;������������h�z�znGJ����:�����\xK�;1���x�� 	ppq�'o`Ԣ|�&���EY��i[[9���1M6�]u���ч=�g�.�ca"�ׯ|�\}}�0��Bgĺ+��Fy��_Eou���p�dFټB7m��'�[��f��Z~a
���dٻk�m��Ӆ�NK2q���U昒���&��ŭ�&�|�I��l$+�.o��-�E���՚Ư�`/$��c�g�O�Qh
 �1�ϟ>}u��벸t�S9u��}r 	��p���Bd	�
�����	6NN�\L�e���"�ɐ Rf'%��o��CS�F�G�ъQ�~j[�}�=������}}�A�#T@�ƺ�ţ�)>�����]�IVV��e&�l���ƥ��d".�M�䳶4���::�U�9��Չ��=��@2�C-�x�����
�'ש�vM�o��P����Fzj�Ed�����e�����]����f)ɝ>+ީ��t���\lZe�9������)|6G�v��+�ԃS�QR�(����}���A�gNd�;j:'c���Y��A��2F�O�̔�$��LЖ�mﯱ���	�0EEE��A��y畭mmu=)���{���}���62h5حSt�ud��|,�͛7SY��uK=)�ou�V'�i�޽;H`����y����W�x��"�w�ճ�����>��Lѫt�vPΝ�"j�]���2&�&�q��@i��� 
o��g��?��(M͉͢������͢���/_�|�B���	�]�^19�y�����4�`���[5��%��i��?X���@/�3��P)�xZ���BEsK��F����I��M������C��k��*�F�W�����JӴ3���e�Ӛ�N�C���qDA�㐮�؝�Q>���.=�Y��g�>.�j��Уq ~~Xo�H������q��jLJ�^v���
�+��*S�����1� ��ݽ8���0vWW-�Ľi�bx�W�5*�g:��a�;��kԌ��Tb����W��{�&1���[hg��Jto�v6@���9r_�ހ�(�L�@ǣ!��y����c9�-��~��Š�x-#0�^��O���r�h���؎��i��۫㥄�ǇG�����]6�%���&��cfo5�wx�3�ގZs,F��ŉB�M�o�,�<~ă���y���L�!����<�e;�B�%�ܵJ��0GWBAFF"^��M�M�����=�a����]�[���ښG��'�}(�_4\�}-�2N�6�ۮB��^�`�V�؋:C���5�oT.����uzNpu���>����W)�&������Z��6���Ȉ�,(�;K�b������ӝD.#��D��[�B�����y�u�ρ�2�2���U^,0(h�<Q=�!ǯ��WdL����LK߱�w��C a����UW]��ᎇ�*W�&kQb*���T�aXZ6�Zf���RS�/u�,l�v��7�c�PT_��y�&��+��!T�ɑ9�گ�m���d'�|��} D4��a9���U��-\}8T}ިy��R.�����:�o�3�.R���D�xb��ܤ�,����K�r��n�Y��'������Eɐ�Ȳkda�ǰ��Ͳ��HK ��( ��߆�������..����fd�?[#o7�٫�ϟ?���5~��MZ���z�:��.Q�]E�������'�I�;]�c�p����e�ZЈ	�&1*�p�V�BL�'������\wnrsߨw5�w�qe�q�֏�%g��2��ٱ���B���ܒD ��0��K>}����7 ��iׅm]z^@ � ~��ugASi�ּ`�r�y�A�����f3�_
:dh)��ED�f>�����!9�Ti�Zi�Vb���z.�&<������Z�_�X�JJ�����I;8�ZuM?�\ʞهS��V�}�U�Cs�/�n� 2�%Ooɫތ��@�O�n)1�4 /������м��x�d&-�׏��v��8�0}R1ᥠD�a���|��!���|�ܗ:[�ٷ��G���W�*M��R�(ޗ7�Z��;>T�)w��]dY�w C��dDS�����#77��P��CȞ���	p�&I�^5�2}�� �e��+�)�L�!m���z٪��{��F�g��ŕ@E>�4[��O�������ʬ�W	;�eꜪ�	�h_Ʉ[E�Iu_����)���N�[OV@
_�v#NM�J��S3��Qii�y��ͦ�� ��6�����棹F�?C**D"�{�Y�#���(�k�I���ol!�� Zԝ��׏�6�g-��J����f��ю�h�W��k��%���*'�N��~VUy�^l�@Ӟ�U��ԝ&��e2��O��=I�Q~�&��t��uQ"�$YBTT���QL� -�kT�~��"2�(�$���C��y���:���>�[������̞jood�q��N����U����kA ��2� n�D\���Yuˈ���M��9���C��"����ހ�7*���(��D(��U�ײ8����%���@<IC>C��g'`�)��N�V��kVڗ���m���������̦v�t��8:�GV�r��Y�퐑����c=!��%w~G\��>c؀ê]��}~��
8ɡߔg��鰤��j���t��LVK�"�c[6r�u�̑��n�G�*\5��> �o����{����?�y"�BB�ǟ�>�`�efj���ͮ>���i��6��P#R�? �C�⬽���v���,[���U����beˆο�f���F!�uh5�?�l��1��5O>�T�/���̓̕<�@�uo�Ʋ���!)��U~�W�@����:��	�l�5�҆��>H�S]A�������2���z1cJݶ�2ǌ']ҪȀ���ܰ�����D�I�A�߆�����ۚ�tX~�}��@Ff�\���׾-�G��:v�Uo	�i�Ϥ-�m*�j��1*C�����ϟ?���J�u�pg�#}p^��2��X�Mv�k�n{��D?��Y
�w���|yyy��6�v�9�k�Z�ga��w�!�P�/.)�KU����X}H:k��_a�}Vd�*�L.JЎ>�������|�ʃ��~ �ę��dz�ؽ��,'��o=f*�}�`�^aDb_���3B/�������J��������w��nU�1G��/�Q9�^Ѝ�f�(4,�M:��DT¾ԇ9=��Y�~l���t^5�0������^�*��̑�/(�l=т�}X(BK ������ܶ� V�h�i���#n�����ː�b��,w�j/jd�I������B�b�id���a
��Z���/D���B&�yxO6��T��-�&/�/�P��\����\� �ꋃ"�P�mX�!������wP�r]�K�_�A[;׀_���ͧG��([h����۫1i��VF__h&COkV��S�4�I�'䝏�;�4F�9��{j<`.w�c.W�l����2��꾗WUꓭ�дM���>��aS���y���"*a��Y �$� �0�s�(��P.2<7�Yf6��Z���A�B�u�`�� ��{���		��'9�aI��Oc�wkQ��C�'c�D���wK���K)O���-J�=�0ntg����~p=|�A�ٳg,Wn��1�o�[��l�8?���^2��X��1������!!�N��oL�
^�4|9�š�ݽ�7q��V�x�T
jq��z��"oL�a�;o���;Pג��3!�����	Z~ni�n��J�y:��ɛ˄mY��w��6����ύɔ_0j*��e|{�}$�H�����:yA�\��-'�c�!ó���a��0�"X�A�J�O�O��R+kiηGf�D�l���A	��o����Q*�
��ܷl8�냎>A����B��������S'�;�����=>�.j���b1u+����S�������v�;������Ѧ��T�χ�Bo204s?$j�H?�%��=>F�Y���u��{6n}Gj~Y#�iu8���]C��|��SYJ��º��7��6�����Gq95����u��#C�v3��׮R�֔�ͶY��O�+T��|u7^��&N]���n��d(��j+���'J6����`�r+#��:�E�Zq!��Q�V�g�ާ)��iRD��y?��� >�	
ʯ�#�ޢ���Ϋ@Ԩ�����7d4�<�R3C�9����_"��bQ&&�N��?����8x���<��w�-�ݻ��2������#���K���k��+�Nc�%��� ��z��x������>�~�AH����a�"���
Ua���)����z��o?=�Q��$fk��e�I����� p
�w^�t��zF���
)��70����It��#b����Qp�(~��eZ�Sdd��+ҍ^w��{����R*bq���n��F6Uk�ĄSw����[Y�a�b'�=g���S1b]��2���%�G��iU��D�����&ɿlAY>PQ�2aW}q~���/��W�p�k��%ϋ����7v��c�!�1����HЧ��°$***���)|�����s�<��.wbߤ#F�4l�~���O����}+{hO���R�4d����S��JW{��f9���F�C7S��֓(S��	$]h�g�pbY-��̽� ����(��Yv��`�#�ƶS�]��8Nk8'Ň��<�jCN2�UJ�G�}�W|s���4656�6[�\+��/wL)ǰ�
��׸����`�"R�7L���e��ߘ��C��n��c������4�L;�����Ŋo���N�܏�����@!�"����F�ۉ�����&b�����L�.ΚȅX����F|)hgkO��cʼ�²'3�u!:/��}���F�pFF�BR�Z�$11���j�Љ<c\T��Λ/�5�"�]	hi�s��^3��{>��Y��@#��<۬���l3�yͦb+//�����̂��bg�ʍ������N}�ng҉��R�3�ja&��ڗV �DX���"%���{�_p��ORe5�lӊW�����U��2ֻ�g�6�����8����&�B]��:^�;rßС����M8I�sBK�ͭX-b��
����-�/�Q���,[;ZL��5 �Z8�W��24���q�p>T���:����j~W�6�D��^z�,����(��!�
��w��_v^����Α�� ���Z�ѫ�o��g?���ЈrT�a
Կ���P&ψ��u���L�\��Д���-���=���r���mt�EGGG�^�����	Ma7p��+<,?��o����$�L-�N�b�<u�(�崒_�ȵ�"�����..��߯�FgQˆ��}�d��L���W%//��8T�y���(��]��^� )3����Z�ҒU�p
�?K�|uA�a�]�9���`e,Z�%���Dpa�EV.���A96�b�,H��t�B�����ǻ�_�*�Y�C��=�R�.��z)�q`Ψ���t��+�i����g�9r�~���,���u�&.	���Y���k{"%�;�t�E<�z�d&k�n�!��FR}�D���0�����O"�4���Fzؐ�@�p���pڿ�ڜ�����s,C1'�7!���q
5�bk�
�0>�����{��3^��.�B^.�O���F-�x�kEl�dW��U���<>�50C7��s{�
1�Q\FD�����4(}���؈���
"���Iiw�Z�X411��=t���X�����U�M�$��v`38����~��aIC+�
�_�i�O�wr�r�D�&{<2?�ۗN$.&�����1�_m7A�C�ݠ���R��q6??����E��V����Ld�\�շ�v:z�����jEt�>ɽz�-v���Ѻ/������������M1�\�cZq��_1�Ǹ)=�6���U!ȣ�p��S]NC��q�n��6�½v횘��H�#ʋ��L���&�eZ�E3�w���Ӿ�&�͟?rd����<~L�b��ȴR��v��N��0R��>Y�P�������=�[�$�,�~�_��1#t��AC焴��\?"���s�Uc��媂�}��������'�ܵ���Z)))iT�p�Uθ#@�gk6L���2�z�I���e�����1>>���y��pm�h7[�N�j%R�0Y���%�$�1,����Kg���zח/�"Տ��#��Q`�N��S��S��Q^
�*n[�ӂ�Ν�o�����q͍�� ��:��������(��,�t��"k���o��D��jٹf7K+�g�h�=�v��O�kZ��=N�7J�֖S���1�R@~Ktp����,����kUy!n��ӗn�-�^R��(�2�gԭ�Qs�U�LEZ�+a-�t�f1��^��V�bb�����P�x�^�qI'hw��Y���8�o��Hj�H�ه&�t��º��%<�X
��޿�Eֳ~}��\�<:�x#}@I���iZ��]��ig\�� &����A\�@�$>� �O%����'����o�/Og��B�π�aV}���;	]�Raɟm�_�i��;���d���gM'ʝ�+{�
7⥠%���D�8jg�en��		in��a��N�Aj�T#��	���u�!5k,�/_���1�Zؿ�)f��^�����(��^�zdt��7���=?u-|̈}���Eq�i�X������9L\�7�䱊IL�3�d�>N��w|����`�R@�5��'�k���� 3N����2�!�*È}C��%o[d �H�d��^�u֝�m�J�=����w�q�?4����=Cd�v�rm;Gu0�����d��	���:�&&�̪u�&vΐ��4��8(�]�
�z\�#/��ppl̋��O8��C?��n~���su��ի��� �7:����Z?o�t�g(������7a�zLmF��m�b���W���bɏ�i���'|���ʩ����O��j�X5���Ѹb@o8�>�M�a�) ��	N�]��K��)����T����`��sGL��h*21A=�eF,,��bV�-�	��������k�>��Fn��!^�;Y�w�=�L��W��>O�LMxUbRY��˺��T,�����"�h{{{�648s�nļr2�XlL�ߡ�*��*BL_�]��J��(��U2����*7��eB�neee.�q=�D�Oc�����8ܝ��0�Wg��9;��RBV�~�	����N�@�2ݽ��p����, �|����u��}vЀ
�3$���������A�_�?7��ν��㹽�˱�����"��a�Q(M#H�/42?�h��\%Đ�_�#D���4^�D��H��R�|��v����)�#�H�L�j���.u���J�ve`�~+i�=f���������}����f�N�6����c�5���p�EO�8ר�Y�1+�	��?U��$b8�K�M"/M-��C���lO�S�#�Yn���*u*x/�K�b)�4��5��v�3��1��i�q��U�����D'�MTP��Wq����A	����yqo¯��#�ۛU��+����1$]����Y/u���)[4��(E�g���.`�Sz�<�c5�fu9�p�}���K��g}z��?bJ�T�泺j�D%OH0��A����d�u��1��\��L�-��{�;Nh�H�����0u:E��ڦ��&7w�m�/s��yt8���vk#8I��%4���(�S����a27?/$�ɦQd9b�a.q�o�A�嘮��`�^�g�1!�%|�ho'�/*g�DPA�ߢn�fE�m����WkXQ�eg�S l>+�i.�՜�z<M�+�q����-�.P��b��^ߛ�E\���U�ư��U<$jx��|P��xt�9c��͈;(�����^�H	F2�2�J���]�ԅ�u�~w����I��\VM:'/��>(��$aQ�"���0�Ў/�%�~p�>2��UpS�BYH���@C��`cklg�:?ٸ���=�N�K�
^�� (I,_-��W/����H3�De|���)UTlE�ʐ๯'�>hU�Ƃ��A@M���r�����!�o����L��[��36�ܥ��2kr5��gI��+,(`�) �&��1ύ!}�����G����x���DDI%�Y��XIp_�۫^_>���!����PQQ�.:����q�k&�7w��� �:1���ټ�|�>gcm��(�AQ��1Tz�seǷ|�h�1�w�cmW�d�o�mhH�����ؾ�Gcr��a�[�#�4�M�Ws2O����:<��a�!M�wq�HQjT�nի�}���QM�.��
�� }��=t��e�]y�Hu��?�_
�E1O.;c;xW������]�����:�<?����P���b���z������b��2g��h%�Iσ��aPHE�2��	���8u�a��p��\N��>���b(�����U�gV*��Gƙ4���1��w���δ��Ï8�ܿ���0wm[��"%o��r�kw"D��AS555�5_�cP����6F)�Tq��hQ���4�ݬq����0�o�� �>Rߋ�{ְx)O���
��.���g	Zl���	׿�dF�XT�@��%�f��Q"���J#�f �o֟�cZ�u&�d�,�(--}�߂�G�!���231i[�(���g��A|�-�H&X� �b|dŅ�vgz�s2���������vJ	�4u��9!@���	�}�Nk��#ST��W|7�d��
-�-�UI"I�.��kE�[�@��Pװ�P�a!�Ǒ���j���D�2�<º�PiM�u��%�'�����������Κ�ࡲ��^�o��D0���+Ydh���y�ԄU=>o���Ğʠ"��7��&�$�XAKkTH}��p<��yT�o7i�n�t������˨	р���R�2���_+�2�m�Y���	�$��rKU�b	�Z�ؚ��rض�wj��l4*tۧD��RJ�g�����lUp ;FFƎK�.�ʆ���c ��cH�i���!�_�cε|R�Z�,b���W��#���VO�z'5�2k������O*��u�lk	�V�..%�w��,ޤgCO!�{R�2W/�ّ�˫�6���B�FI3B3�g������W0:$_��M��y��K'�=dқL؁)999ݡ�R���~x��=¹���@ۓ�t���Y�j���x��)�~�y�y���K�45|��y/4;/�=���qԌ�%����X�D"^��]q~�����S�eP�b`dڛ< [4��繳��+G	SÁ�����]�����Ɯ�w��uW./Qe���-�I5�Jp��3���\,su�%��d��!d\���cc!�6�׋x��W`4K\�4��P�toZ�t�%�kP��/V�ݐ&x�B��h��L�Ϝl{�=R�!���p|eY���|�Η�ߘ��{�Y(�.d5Hۇ&&?b��XZ�?�U��i�fU޻���7��������fg,aj`'��Dp��ۀ�L#�ֿg��S���,Q��|�)\�ztsbć���V��B8=6��P:���b��r1o"ش���4#>%$����O��e�䤽��b���c��5S��/���Ke.����##&�q� ��ā"� *�Aȩ���K#�[�R�H��*�B疸l%������q�����D(د}���-�c:����� ���0#_�Z)sR�|����^r���Ћʟ?���ߺ5�A��P�.>���@Rӛ�9�d�dĀ�}z��h���AV��/��������-��n-&z�ۍ�P��Z �_�SSt\\���.2॰)�v�A*�,�V�uz�%1v~~а���s��Sx'4�"�Ǧ�0uJ_a
		+aY���FU�z=��ʕ�**D��˝��3�I��� u	@�Z�(���T��k����]�v�a�$���C��7����FCI�[}�YGb4x*�s�dT�� �u���������mBX3�d���DGG�ϓ���Ὣcy_��\�;-���k>����UJz11;;;��x�--5�>@��ІpݑR���r�]�[�~�8�����,��5�K��r�"B��	0<��"�B���5���MQ::ԧO���T�+��<�Um���U�;�Ძ[Zd�]�d\�o�g����iA��e�}��WQ���/ �vM]z���y� ���TZ<
^�r'iE����MA���%%E�E.ꢺ7�уV޼{w?b~���v���
%���Ce+o�N�-:	ח�hd�9�j����S��<iJ��8(��]kWn6Zp�*��]aQ���ȃ3�味�;o��D%>�-�~��?�yoC
��]��K�z@)d�s�O%�����ӏ'�$���5��_p��{�(� {� y����sh�V�����CA�������Ϸ��cY�/����T�̊��R��Z"[�11g!�*�QwM����[J�OWy�+���6��ʪ���ٷ֠��y|:,�G���d5]A/��+�k�u��{m� Q�� q汎9:�
:Ӯ||=>�S���Wxf!d.���D�LA�v%���g+��Q�Q�ϼc���w�2Ӎ؍t�|||~�Q��w/å�eQ��Ϊ�����C��� '��4�H[�fI���!�`�S�R�׼�~?��ȸv�}��-��MߟD���
d�d:�_����w��_�dM��d��C��uV�vXLT"�P��"ۏ����H@���&6G8\�Є F&�G���p���҆B0��].���vm�O���2$�}g����;
�<<�?<�H�N� *���*xii�>ɠ#!�+�t�aV?��֖��./��q椥���566�2����\�,�`�oQ"����	�ȺH���%�S���ttLL8�6Z�m���Y��-�����	Z��x����eP�M�ח���^(i��1!���Pa���%�E�N����U9��۷��������\e�W��n�H+D��V}��e�3@��P��f��'�{)��h��~d�ɺ���O^���_�$��"8*ZZ2���p�����/ց�Ti� ���\���	�H���pt����׍|�/ (Hy/N=K�u���^�!%ePw��@g�E|��eta���2*\�:����Y�*4
w^*�#c��]��#ܐ?j���'!���H��x� 
^3d�\R��-.��h�`0�(�Iz���H>��h��[��Nv��?�������U���/�H(�JHUeB��,[��ӕ=3�AvO[6LE4�$��m��|֊AѤ�4��ÁNi���xKRsj�!�@u�/�{���/��WT���S��Sb�``�e��O�?����U���0߹�h�B��C�ލ��=�L�-�����.���^�b��|�3>$֌P�����}2b�P�ŭ�?VT��$Ň���}r/�0V�HI)/_���ּ�8*,��`@��Ŕ�����ë⧧s�Z��d[Z[���N�˯w�P��L^$��'�7sȄ5l��?#F���Gfg����������F�T�/� )�c�M��*� I��?��0O
��&C]�1АU��6���M�nrp�f.J}c�8W�z��~���ph�*	�[󤺎N0�ӫ182�L駔�0_�Kb_�@�>��E�]!�Ȝ�D���F�F��
U�����ĝm��A�wCe����������p�<��i��B�uF,D���))3J8���C��6�#��*zC8�-K��t'�2Ι333c�Z�$Nr�_ӯ�d��9?�m���?f�H��:?v8!)���#?g*���/�s���:Exa�z��-Φ��U�s*J�fH�Wf���\%x�L;#'ӡ"pHLL<r��֢�C�{*�u��w_d� ���+[�p1��>�o[9�6J�@�IJ�C۟�b
��d��0����������.�Sd�$����Қ]x���Drد�n���"��w��NՂ^�7~6pd�H�M��r�+�f����Y��99o����� c��($�����d;��A�����w�B�ņ�^���ϕ��c�C�.�	9��-��wf
^ܟ'�|/��������~n��12r1�k�d�U�b0<<"��1�u�B)"1q��"��.R3hׅ�Ƨ�\I��>�Du�(D&_6� �z����q	O�6׷H����׍��&�$&^��:7h����E�9�J^J�xi�R@��V���Z�g8�ȍ ��T��Lee�Os���6Vۋ��<9����d�_������HZ�&g�����c��pW}��1-�A�'�n�E?�W�esJ�Tm���3��=�����<����zx�L3��k^���;��q��mx�"+������?�,���~�gJ�e�p�t}:�)0JؑY����L�[��=W\� �o޼%��_渲��Le ]���h!���"
��������mΣ΍�pⷤz�2��>@[�D)��6[�D�S��3��l#� [����WT��|�����#�T�/���
ߤ�"pE��~�R�$wQ�@��b�PL\��	��x/Bз/�8���ܸ��:^�qیڼge/�3��@�|�0\�;P#G��4���@M����#9����9U���g�͇�#[��!|��k;;.�{��.t�#�o�#�;�����GF�/�e��&Ë�YTc�w�Ѻr�}����3ԡ��ݻ���g���K�E��}�ާe����cd�����WG>cHEQ_�u�xw����{����8!{^g9䮑�f�ՙ�|�߷�/_\ʈ�s�qI�YaT�u5J�� ���c���@��Ј�U�h -kR@@MU���FϲC�5,D�����l�?��]�Lp�' �l�W�ɕ���D���!�� ����No�;;��)��N��2��7��sUS�ګ�����������W��qd�{~ve03�\lYn�EX��H+B��e�Ydw�������B<O����tEq�J���ش�����6
��E55�wz�::T�� e��� m���"B�����t:�����-~~PBe�I}CJNNE�h�����Y{p��&�;
�n�Nk�����&d#�S��2*�F3ȊMR'���� V|.8"W9�"��t�������v��4'16P��'�<UE�'�ϼ���k��G��4�ܮ��>!Mֱ�X9Ę�/�JgQ�J{��ҀCH��-�|?Z��Rm�'L00b����׏~�E�wt�BW��״.�s��Ǯ��\w��KJ�7���Ҙ�����"ڲ뉔����"�����\9�J��58��`.��P?������/m~�Y�Ιn���Sމ��K��KE�<&,B��<*Hӫt��������ř�����9�d䠘5�]��5����]�~�ODu�T�@�����o��T�0���L�ߘ��7��J�*w\��S��܋]�����\��1t\ả���B}o]��ռRaW#gA�������g2ۑ~�vuF^���74 ���P����������/�u�e�(��01���e~Oh�wf����pk�7/PLԞ��G��(
	~��u��PtI�(���6
�z}�@�D�/a�o��~�_���׾�3�uXܱs���)j��!f��A���r"Dd�ȅ�#��]�%��}}}���F��ύ�b��������N�_���(+�(*fm�xn�"����ڼR��Q��5���d1qq}}}����1�������������I��w��ƖOX���N�0�y��,`��"R�M������V�
$2��	'�(Yiy�����PK   ���X�Qw�M  �M  /   images/4a2284cc-1baa-40d9-9462-4dabdb252300.png )@ֿ�PNG

   IHDR   d   L   �   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  MIDATx���`���6|i�aɒ��؎���
a�6���R�@)���g˦-}��/e��=Ca$d/�#�{kX���Ϲeg@hy�����Kz��g^��C�.��RU�I�L�SG#�$8��� �bV��@�d�T�D
F�c�Q��+����:Js��ē�'��Q���}j�ܡC(�D��F��������j!�H�'�RHE�
�^?=3�w,]1�4�'��-HŴjJ�O��(�r���4*t���G�����o])==EB4��j��jP]���#��z���,EĖIR�}Z"��	x<^X����S1ѩ��)P"�4q� ��M�z�^
z�@�
U�/�q�,W��.�V�$�y��=?��R�z�r���ӏx 
u(�4j3-A��1��VJ�9f1v,�l�
ni��O����S�Yj@B/>ġAB��<MDF��I���Y�e�4��t��2�ڥ��J�C~j[&������Hng���s=�s�D۪%$�Ӈ��Fd�z���O���TB��b�j+
�J�Nw>&<A�<��r̆��Ŝ�t������R��Ü��0[�J��)-�C�Q�$}ua$#`�u$��
h�����r��:�I�"��`�T*�B!Ҽ$tZ�;�pCP��(�h�� �AK�e2bd(��[�VK�K���J���D�H&X��
����4\K�ƨ�եU��k8���p�w���b���P�P0(���X<��3ψr�.L�L&��~����2TP{���䶙<�d2�P8�B�1�1�Uy�������gQ��Ci?���Q�G[���ଢ������r{$_C2��RMiDuP
�OA5N�#�)� џ�ծ�4{�3�I9��RK�4�\����Z���x|^�ڽ[�7j��;��ˉ�G,%3����;��p���
�)7Z[Z�x�b�u�̞vA�E��q�vTQ���B�L����˖.%�&E羽���������E��=X0w6d��Z�H���t�`)=#�*����Z-���B�]��3�lz{1�t����wQ?s2�t视����$-Z��pͻw���
�~��:؎�I��M	�a20B�� M �TJ�����u�Vl�R���Q(IM�+@k��	?lF-fUX�s�zE�j��)$+?�s#AY�I��J�	T���F��d�
��`6鑌G�����*b���j�j�*k�2s��A�����(/-B�*$��{z��>F�[`2h�YM���TW@.W�z�:5�6u�{4<�'�[�:� 9=� ��		��~*E�&��ڎ�0߁���)���
j�����������3	����Z��jR4�iuC<S��M,I���:\8K���n|�[D*FNQ�B,%EPjEl��Ԙ�LFvU���I���K��S���݅��wDY��?����!I��%�\(�/��d6I��$��
�R��v=�?�1�Cc���9��M$H#�d>l
x�YS�d&tdv\�I�Cj��[")�!��@�P�C��
š�z�Ĵ	�:�."�T�Fݣ�Rƌ�Ø��x,�P$e��ꗡ'��,\_��C�%���IY�)2C��縟z��ԯ	�<[.��>��&�ǐ�;�Gm'�����[B�D���:������zz�!%a�ۗ�}�e(��
F�H;�j�	)d
I75�P�Tb2�"۝���?��0�D�vR6=ia~YÄL@̑kd���"���F�r�D�����i��=ߢG�C��/|S	�+���L���#���2#��=��s�P@�ojv�z���Ʈ=�$�)T����o�$�WV/JQh�f��Q�C��gv�3�X
y,9���_T��l��Q?�	�}���ns�~��D�F�ly�����;�l��"��6'-�]�,(U�o�$���8�j�@��a�EN}�k�NAIr1�O�PA� �I�Ԓ����#�$�z�Y�]�3��H@�hK��%��^�0����3����rL�`��c�~�9*�c�HVX��������q��ᩘR�y$O�o�cYV�0�0�bq�p�P��0R�թ�8��#8�3�=SvY�͕j�v�v�_�E��^"�C��c��3����AbF�m_�ŕ^������0��Z,���=ii*Wc�Fp������6Kg�G����p{"_��\Y�J�	���<�G�:�6�ɾ�$��b9�X|:�*��l]�����c��0�� [����X�W(	��o���բ�c�d��?r�.W@��Ң,�w�FɶkPZhA�>��h���阆q#�&[���nV�S����3'��}��7��m�qϾҜpvU�����둟|�z�3�Q�qĖ��'-������X����y����?���/��|v��g[ƾ�q���l�%�_����6�]���^rFE�׏���gg��'�%I������#�'i?��s���~���[>?��}�+bI9�N������o\p�+Wl�:��wuÞ_��Q��c_��x&�y�+�o]w��sN:����m}����N�T߶x�9���y���XU���s�|�U����|�eu-�[`�rؿ�3�2�ӱ��Ks�u-K.�F�3!��(��8}�a^MN{r�M8��@#���`G��1"�Cd�#�`L�	9����	�d�BI%�������)Pi���MS��F�I��)��$��nۥD�x(�F�G��uݱ��wl���eO�^�@�ר��Tx����Ɉ:���.K�}��x��Z�h�uԱ��g\24��L���g�D�:.�8a�}��?���2�uX�W�S�CZtz�L�mX��&�����I��lrڪ��d���YV'��j��2�4��a�{�Z��s����g¾�w;�>�7eTy��{]����S?5h�X�����'�&���0�3��^�i�p@�,�xz�����������<Ð�ɰQ�XW�?,>j"�NAa�v�":�(*��$9o79vb$�mˈ�]�AX5

���8%�V���S��`M:��p�%g�w�%�y_9�h�^�� ��oF�N>.\��P6�Ci��ΊB���P*ӐÍ㥖�0  ��n���:Μ��W�ӯ����j#	�x�q�)Kf�a3�ӻ&��;��y%"��tlɒx2�`<��6Eפ��0=7#�����"릑���q���/M���{�5|Q���z?Ci�ݮ��5}%E��$�%ɷƓ�4�W�^����zү�~�E�r�AJ��j:5N���b$��Aѽ�ϧ^k�IӚ��]��Y,F��$?.%���6�$Q�~l#
��		i5J
#�)���(\6KI��9{���	�C^r�	� Id�~
�-Q���0�V�Ӗ��W=a�j	�X�R������A��	�$%�V58�!W{����"����wQU�L�9��#i�����d�'�{v�E�aƼ.��`B2��8�������b�a��X"̷$5�y��tYQ]����"B��@��j��⌺8�v������C3���wN�z΂�������A�Pa�tOӱ �S���X����>�47���!�s$5�%��a��q�ԍ�ՇZR���R\�.٨�2r��~#�k��e9�)=�o� �P�O
�y�w7�C)�#㴄D0�u�K�`�"EP���ɳ�hwbs�-�O� �5i��>��R�ڢ �J�,R/J�K*�󥢲�i��ȯ�L���eȜ��0MA�YCR�e��uM��V"��� �h�(F���<�F�6b�hK�ꧏ`Gw���ťu-xb�RS�h2#r|kq��8��2�dX���>t��"�22*1���{r�͹ｮ�%C�좚}-�(^m������O)����p~Ó�ՅF�uSï7�U	\�мc4�s����`iN`y����%K�]V�Ye����D��}��9�P���--���zʬ��w�j���w:+����W�nk"�ռ�VSQowFW��o�0�?���<�5������m�0�ϫn�>�7��Q�Gh�D�h�ǽ�K�=���LM�MN���<��{K��V���4kuE�DU�d=��SJ.���H���)��39����ɲ���M#�l¢��"GV�tZ�O��p�é`��_"�p�dFm�;�u���"�(�*��eG[q�y'IJ8M"U@� �<8{I&�fVGpl���7��ɫ�n}�פ��^>����ںs<�%�����xx�=�ׇD�SVu=Ų���\�C�%}l庳���p�	�c�F6?p�C�����&���gTv�Ub������Rl�r?x�C'<���O���股�n������>�֘}u�ޟv{͕;��.���·V�q��a��Ԟ����f����ģ��[���+~FN���y#_�}�#����QuvU�-fU�K����?F�9��n~�s2�"b���^���=�>�G �|���ls,�1�x�����]�x��6Ni
������׌}�=Q��qL�9s��b'(�]�>��!9/l("�H
s@D���mX��8�|R�C�7����(����|�������[Fss��q�ܿA��VV�����펝c�Y4(|�]~��f��M�/?9�#BA��(:�ƻ����`au=���Y���6��A�f�p���3J;�f|�Wr^��w/!4ce�zr�W�i�Q=4�Y����!4T�r���ϑ��ˮ{�쵄~r�?_����uQ�/��>Ee��Ԧ'�ɥz���r�G㼤��{��6�k�8	l9����N��dɆ~{�����g[r�h��֬ʿܭ΅3����I��ءK��?$8NJ�	�����4B�8X����*N�K�D#I�<�t��"A�Ŕ�V��ۚO���8��H�=[���"HA\qo��]�+0#c	y�롂"��^"�TT%Y?P4w��K�=j�LD��C���z��d�#qE�� �[��Sٍ��9��BX��zf���$-�R��\�`o���4u���T1P4o`��p�.�b�,���D����G�Me4)]0�a�]��f�ТWD-9�z��D	�8#�ǒ�g��\<�v�S��o�pCjfϞ�D"~�qHM0w]zT�P�����7m[�7��KM����L���z4����5��9�N�˷|�W���ګ?�4{�|n��߱ɺn��[�|�#H���QYO;��G�&?L�w�j����]�o/4�CW��{Ӗ���I����۸�1��M�Oc�T�L�xf��+�捌�?��v�����T]3w�[d�=�{ޣ$��_��}3i�q�;�T
[N*�{�ﭵ��@d�j��?P�6o�0{��������?{m_�"z��<�ě��{��ͻI;˞�=�R2��gT�ݵa����Pz�ܝk,�ྎ����`)��@�ÄP��;va�$��'&����+r�L���"�p&x�˝�]�G}��7
���M
Ņ���̞
FAMe�MQ�^�2�*(�׆����!s8\os��8����g2�#�,[u�x*IR������=�265'����2�g�ԑ>���\'��#�H�\\��tUfM6��q.k׆:��M���C�:şI;��M�'M>$Yd�P�X3ݦw6��+ca�cUGz�LNq���,��i���m���fo3}����`;�]�hS�Y'�x+!Y��1+C�TLd�y�g=
�(A�~ELa.p9��F��uV��AL
��.��O���;�0kV-}�¦o���t1B�<R����<�dRߓw��,���/0�$⁤���|g��127�76�ܦ	�|ۘCt�o��>��L��E4�]�v�{j��6�|Ȍ���7�>|�4�y�����ɡ����.�����0Җw�L���S�L�w�E��l?�w�m8�S*�>j���r�c'i���X�{Fb��	Φr[H�1Hm��T���ȑ�L��������Im������=v��ʚ��u�e�
�����>�v���d���������~�E�F�쮂
E�aX�!,��G�s�ar\��k(Ԉ�MZ#3XQ�Ё�7y�
Ŝ8 "���ц�E��X��5H�\J�0@ I��kLc�����#$�F�
�ܔL�V!��i�6��SE�|Q%�&iM�ѓ��ȉ�eٚp�>H�,XTO�5R�t�Mmh�|��4A�mRy����M��8mD>FI�J�g��,"�h���-i����3mꂢ� 1����?
�4�&M����T�L>XB�$M�H"!��D�$�e��3����8�|�����`���^��7��U�{`�fc�<�r�Uq�T(�\q,�L�H��\}'&=�xf�"���I;7s�;�_��?�KR�sˢ�����t��$w���{�Ytף����t�%���?����}|J#�ٳ�~䧽�gP�{Ϩ��꡻\��;��B���s��A����#�z�җ���I�Rݗ�_����'���'/_�D1���%[O#m,�z^8�`�����^z��w|�nZ��`��'����OO�Mb��'}���}�.#?�_gVv~v�MO�����ڱ}<��|ڕ�|/i�GU���W?����>G�p���^�a�7��ƹ�ΰ�x�M'� �'������=O�v�������Z˒j�w��_�N�?l6́ݤ�NҒ6w������z�^z���VD���!BEє�u��x����s�ϟ����dJ�"&���J�<�*2M��zo����fFAd��&�֌�� t��̳�=�1i�#$B#'Q0U@R.`�+���P�j�Gu�3O��15�>o˹�4�'�UZb|��U��Z�h�PѲ'?[yO��d�ϟ�_KDc�Ŧ&���D����U=�7HI��n�s�?g��R���������g	L\ʾ�\N.f=�����^���8�zb㑿�2�ؤ`���'����*y�_=�>i.������Q���Ob"��1@<�$��B�KC�a*�Fjڍ<(r��	.=�c1��2ʋ)�'���O����O=�T�~��"�8�S���*��J�8�FQv٦���9� �Ŷ�4N=L����=I�5D8
0�W���'31��|
_�X.�t�TX�~���A���WSI��<�8�4��)S������g��`T�mVm*���&��3�����g}%&Bn�d��6_n�[L&e1�)6������O��ݮ�|
��x%MmR\�>dxʘ&h�&M����0�IqQ-��ڮL���s�a��	i�k�J�:'M�t�m8��J�鬮W����f���r��i�M>�j��>z�<�!Z��Cr��0S��ڵk3ZA׺u�p�EaVUy&#�,��I�$gVt̱��~���\�B�%u-��/Q��y�Q�ٮ�)e=oR`v�����ۛ	¶c�b��f�ۤ�;�/p�?�1A�����	.o"�3E�9)WLP�Ob�rj��LMo�ս�_U璟�_Vײ�4�He����}���(���ɬ�F��=��<r!�X�g�G(��(�S���[\�ڋk[�&��zN 3#3�9��	��U��U�5������e��?"�Q��G���+�w���R�2k���H�cF�W[J!W��Z3�w=�t��/ҫ�^�	��9I&�sif�g\ISt:FGG�����t*��L$�R� �@t^���__��u�wݿ����G���y�*+���6��7�_��o{�T�ą9��P��?�GsL�WF����:��"3�P��j�����u�"҆Z�&X���@�IDﭗ����_���^>��\Ӆ�����M'���R<��������X<�\���;>!:fq��?WWt�CZ|1$q��ͷ����ӯ((%Ȼ�����;�_FqLűE����#O�ʚt�r��}���<O�������5�횰��iM���%���\\k�t�r�?������¥���:��I�Y�r�5�j�ot�&'B������u?�ZZ0�{y&���UK�b��j��7ߌ_|Q���/�v��"[�Ò(*�<b2p(`�����;8����'k~�c�{e�� 	���և{Ȏ����6�f�դ1\�v�F��#eyw��CT�� ��&�9�,� �L^�ſ����k�b3E�q��'o<�ie����%��Ppʃ��Zn���s��w~�[z�Fa�><u+�}=������n}���)�}A�e�}ν�G�ȇX��8Jp����
Lw	��+T�Y��ny�w��(��e�T5�K��)t9���ž/���Z�YD��bș���y�@�_~��,؂��B��Ո�u:��G��K���j��lq�'�Pn�������=[V`��2�X�Aq��# ۝�>��-șJȱ;����')�pV��6y=��ٞ#%MSIg.��,1��qH8�ZI��q=Ԧ�t4��e�A�X�o�^�6s��r�}>���Ӓ� ���xv��!G.'�����L�F6k<9{��t��̩�r�E�2cx��ڔ���r{=J�m��J2�J�8��ˍ@0���΃����M����!��"��TA=$���(�X�4����%�>���{-y�nd2���J�YB;x����M������Ƕ-~���_��]G�j� �E��������[���r�5��cs~�ȶ��"�%��%[�%	\���?_]ѵ� ��O������켏#{*�<E�S�.�vf7�o:��އ����~t�ⷈIFj��d&�}ѝ���~5�ET�9
s�����j�g��[�����-�v��ӟ�=�R�[ɏ���^'����w����g*�&=��&�i��W�7�}t��4����k���	��P0y˱E���s�{g�����:aҙxG�l�i�uɹ�#���cMW��L��B���ބ"���p
�cE�A I���$SK� �+c)#����YKH��ts�����s\db���D@nz�e�����3�,15��:�;)��z^+�I�u�0�����3��l�����6�2m��Y��M��y3m�˪�B���:X����dDxգId���P�/\������6�����d� ��߅�0M�_�!-�"�l�~4��'�Kdf���}q��D����'q���0w9�˛�6aj۾����m��=��78��?�{�U>��_����t�oH����v���_�r��S;\��^���������Kͳ�����X��sb�惜:���Č|Һ���\}n���T�ؿ��s�̾n�ڤ8����-n���>�c��{;�3��D���,<��{��PX�mr���m���^N�֔P�or*��3�`���tڤkz�xfJ6��T��4[�K.#"���T�����9q"HX���QEN~<�O�P@K8mV��7�����nHҒ�3�h�������� I��|Bn�ٛ\�7�Af�t�CM�t� ��4���:���f"����.t��гU��܍��1�Ȫ���i�x,�_D(�9dR�IګُP�$�*���T����d��r�=6M�K}+cb��Y?	��E��'zIc��'H��Q6kt���r��v�_+�:��R��R�o�Lu��%��}�WK��^5�&���c�i%���ȇ����,��Ah�{)v��Ŕ,�MQ��f�( �Q>�Fnv�4t!0���x`g��ǽ��V¨Q��UP`��E�A�&����}��O��2B+��r�'���x��[D����{6��N&\��K���W/����'�Y�����P���	%}���U�����D��׶�Dp���&�����]���7>ID��Բ��x���<�KZ���E��%�V�V���`h�����p���#Sv�9U_T���)o�ա ���g�u�K��]E��^U���ݷ?���;��lp��M���!����<Bm�}챛_$����������9�{zȔ��Y��tb�Bj����<~�}��z����Aˣ���2HҎ������႞`��Eسg���
L�߳f�j1�9>!"�c��.􏸡�v��Z���r�T���E6Z�Đ��>^��q$�$�÷�G���O���z�m*��4Ur�C�|�uԱ��k�uO�wy��7��J^y�W+�g$�˧�m4w����	��K�.�ܡU$Bd~@�,�<x�;4�z��7�6��e�'�-ΰk�{�̇�M#������^�	,�)~A&o5�%1cx�''�J���#y�����֏v��p��,�W!M��q�)*Ϲ��[�'<����P���O];{τ�4S��]�O�Tf�|�RGj��5��-5JI�K-��q!J؈F�i4����S�D]j�!�}p�&3+���VCR1�8b�2�ĦI:)�/O���5��F10=i�f��J��Z�� �Y��-�y�_ΉS9'*�O�X�Ғ	//���{%�ʡPHҟ�����8�	_���ºx"IfT2q���ee,%�S�55�cIG��}8��3��-fc�m~3��&"�8�F����2���e;��������ǽ�f�eN}'S�f�9I����X�/�����V��|�>o�3�J(�$�z��#�d(��(�Ԓ�:��%El�SP`BQ�o���JeJ�!W!e�2�p�g;�"�&��'�
ܷ�v�����Z���%@�<d�x�\N����d&J��f����D�fma�C,r�:�]G��{,�Y%vc�*�C��Ix�F-[Ě��0��$V�S@%��s]<��;�ڵpMe�omk��g��K2�� �4�<�]�'���z���Ⱦ��Z�.��
�X�ƾ2O�1��:*^��F���������ԔXEr(32������J��$1叉��jW����h�nye�!V�� �@���,�ze�V"H���NJd�+Q@D��c$���� N�LNM�U�J*�h�z���)Xr�<�;�ǃc?�L�$�ǉKhf�0J�+Ğ��T �������`H�=��%BE�C���g�H�Bg ��0�:�����!����#�D�)�J�W?&�;o(.��S̤����+9�:��^W|G�!w�[ɇ�1�uB���n����C���	��\Y��guЂ�kB�ԋ_�j��ߋ��j�p��45A����t�h�m��JB��6��\��[P�e���'�E�0��B��p�	��rWt����
���&��R	s|��/��E9İ\NǑ��賐��Wh��uL~ ������� ���
�!ݣAa��K�b���@M��0�mn����لD��ۛ��dZ0�|�Y +��~��Κ*a��01>.�z�9���]�c(G`C.��)���	*�!nJ�XU�#H����?0�MP��Br0�7�����ᨴ⯛R�+E߻��[��:�4�,@�C�I'�"�0�M/���6}
���!ы�ϻzY�'I�9���PG=1'�挻�L���iF�e��iJ"�J�M�KK2{��F���L��a����S��E�;�NՂ��CY$3N���vTq<����6�Z����(��(��g}�mɬL���#�1��C�5�ls��^��ы�0�����{�h�C��O摼8��G����D�q_L0���D�t9�ԕ����~��OΪ���w�a8���l}�=�0\�N����-�P�U��N%����ȩ�u:�kx�$K�EDQ�T�YLw0���r2â������^�"#S�������4&(���޲�(q�)W+Idb��fR�9{z|�/1��f�IcZ[>�1qغ��Y8��ԥB�3{���=��_E�ʠj�dZ2%P$���di
'O�<}ϓ+��M�I��91��{��r�fd��x�Gc�ta�o'�^�g�������������X�CrdtYf̙3&��[���c�.�E/N�G���ӕI��&l�ؤ	�H�m!�B�Qo{��$"��iK"*+�W],@�`���r=��S ��<K���	��d�4��]�1��E|)���G�[5�́���L��W%b�\
�����v�}O��[�����h���p�C���{���Z���#�~���qP���׉���vj%�Q@�ଅ8�^��*��?^q��\gz	��ř>�27�4����\��ib,�%���XƩ��,�00:	���Z��P�.�#��T���9<��Ox�:��Q!9�bz-�o&)В���|���H4���1htF��e_�Pip�ŗ`���o�C����l���`�)���"�� �̘�-�':��&A�iU�ت��M�BR��ih�m�1v�8�}p�<�#�}��b.��EjJ�o�@�*!6�p%	�`I=�c����!�{����g���:����w�)�]]��x6�b���ƚ��z��G@�ވ�(h�%��&�~����Q0BXq����	O����"��A��tQ\Y��ǅ��#���+��5de��.���	��H�r�6�ԇ�ՈҘe�z���x�!a(��D�H==����D�+��"ϟ�@#�0����~�R�}w�dZ�*R�ȼ���O�Hg��w~�|6�pd��h�;�n@�l;�;�I,.0b��H�bih��Cj�	EtK�UNF���$*���d[|�N�3��u�t�*�N��!�9���CMIQeq���(�[��i�((���Yp��?@C�_�d)��Y�y�
t�C�)V�Р7mۃ�v�"W
f|ߵ�Z��"?s�B;�'������rA�Ta�xZ )����21_T��?jȩ�E�n�M�ڪF���q��<�g�(�T$��W
�>�����L#�MiM�5��5ob��g6ȡ�؃,S6�g�ས09A��t���:x�燖gB�(�-+)���I:c�׭�/��Ƹ�&3A�=u���k5���$%�ՐT��-��A�vipL�qЦU��kur�4�M�k�-f�&ƅ�/1�zM��o��,�H���q�MV&�7Fmq÷��?B+P��9Z�������L�O|AO�h�'d�r�����1�Z�=���+JB�]y�<�����b�SkK^^ہ�*䘥8���N~��|�T ��{|�Y'� J���w���I]!�9Q6��
�H��࠲{<>���N=�����G-E�	�Է��0�Ӝ�k(5f�f
&�AU����K_��'�H�.}R>���Y+��� �FR8o6�.Q�/���9����<�ј����(������)V��`�4�/���0Zc"C,���B�d=�C���Fx�^��#Ɩ ۑ�k��t|��77���ok:NĢ8���0�OaC�A�?��IDWD�d��`������v�������,b��g馗=҅�Pnv�$Ȟ��l�F�����
~>ӄ�:E�J�g�Da�[��v�~��]�GPPP���
�CAl�ш�DԅH�e�)�8}6I�;���q���zC$b���l��L:�@u��b�sm+H{UHh�1c��hHˑ�걦)F�P� ��E���͜~'�FE	�Ә,ej
*��Ϗ�_(4�ę_��9 +3����ixzt�|'���S�M�Xv$����i�,(#��!E"��CE� B1�֥y��>t�v��Z����t�5��91)n��*�p���؁��|�N!��o�c��4Č!�*�6��8n��R}�������*J���Ϥ�dߝ>�2#����{\����%Ȍ��P�P��t�{!���q�tF(bӬ�V߳r�����ة頏��2aP �zN;um�B�SW��5y	v�엃������v传�:�N]*��5{�;��bho�p����N ��3Y]>k����T�a0Y(�J��TT��m�]��g���p>T��m9���*��=Q�p�Ho�8>X���G��iS㱯ʰ�ċ돜��5�P�_-¢�(��`G�G�GN�'-�o֔�*.�?��Z�ۮB"�����򥇼?�[?��������c9 �ٗ�ԏ�&��:^�-k��3��!���a^�'3��N�?���1r�Qd���;uN0�}��A�ɹi�	\Y��0�����"�WX:�Ǝn���çL�ӯ:1<����?n�b�H!/�?����hi�p([D_|fK�(FC6�sF�h�r�tYE ��1A��}��������E����"��aL���m@h����V�����O��N��'�u��&��©#��3�"�b���q�� ��h���?lG���wb�Jt�w�)�?�,_0��ѠJêId���2���,�����,U��TA�H۲�'"����\ԡQ2;���b��X���Q�:����&�y6c��a�	��߄��L�m9z��m[�c5���L��/>�mzI���~\݅g��~�n�ϩ �$�c_��K͜����=pM�I�Ĝy:L��!����N}e������o��§�6��WT���4	6��%�"�Q�N6L���l�FYV):���e©��w*L��9�����=:�#ht�z�^�8�/<sHp�2��či\���%��aO�ep^S��m���L�w��Jn��jl��uA��<,-n����I���~B��ŻQ,kp�ʟ]�w���ӖD�8�x&p�
����df�UE�M�}��
�0��KozM��'�q���gN*�v�G�{�q�m�8�(��3���S���>�	���Jd纠#6�{���a���I�\9Ǡ�Py �������[�����\�A!�Ͽ�w|�cGHǒ�@�G�?_�us�M(��^��щ����v�2��=�!�NHt���mbpJ/2���蝠�>�80������;q)^�@�;k@w��,ɔ\{���(>�����'=E�1��X�'�t�T��XJ�m���Wb� ����c��N�}�O�E��z'1�.A*�e���"��=�d���)��C�C;����O4z^N(�^\�g�ۛ��]'�Y]��z��τ����OCJiZ ����d J�Y���E:����PȂt�N]6�a��s��,�F�q� §��Lط{�G��0ڼyh�*��� ܬ���c����g8���ĝ���_��)�����~���ƫ�V&��$?�೐�&D���\�]V�
A�@�<�Α�,����'��C�	7�f����
	1_���}	�ӞL�6���(��4���(�̊̘�HLJ�(�3�UE���9�86���A���+�!�tAN���n�������%G��|���@DbC�������x�����%&�P����R���- ����ށ0~��xF+����[���+O�<�����(�i�@�QAF}HirD<�J��H�/�@�©)�]�C�N6R�\Y��/q`����:����,Wf:2H��D:=}l�,)�X՚fI�Oku�b� G1���Q�#TZꑟTJ��<J����5�pD�!&)@��4�*��0�!	!'��(�l�V2��*Ddy(	}L���<�Rd��`MmED^Ohp!�+��/op�X��¤��|�tP)v����gb�ii��Ł�L�3��"_$��h�40
� ?� ��P����ȩ��ee)���WD��+��>�H/U��0�OHDU8��s�"�3w����??�H���~����(��(��c��xv[9��vX�~�Z�Ɔ=U�✮S�mO
m��������2,�0"��X��ǅ[i 
�aL�#�x�S&�䫡7г��{�W���F�{	H�
	ja��W�Q���RHa^�-n��`��f�(i��f?���l޷���AHkY�N��`��>fCOZ���<�����.)�RX�����2�|QPM�f����f���:8.!����b���D���d+�� ���%�P��7�zn5B}����6s�髦�z�$ӑ�¡�����bj��,e���w������m����� �x'���زs��(��vv��!a� ��v�)�-�FB�'���@���>�!�B�ԼbCS��L�c�{	�(�G�[arì�F� �����Qf��JDXj���	�&��A�u.��Y�ˎ8&#��H(�a^Ɖ���L�����j�=c�j�SJ#�U�8N�}#/웉�Uy��pC�V��Q�@�,(�d�$iX��'23��w�y����{��)Vi�p�J����,\��[/EHv6�s;�dGɦ�sCzB=5�l뢶$����1>���ZFW	��i���b.dJ�t�>C�% @@Y� 1�=1ī��"�l��P1�4�&/s�~��Z��kP��x���&ћ::�P�CI���e�(6�9�iU��f��%�m�;������.;�rh�gs����ޚ�5G�(�/ҋs}?mM#����AG��+�VBWP8��?��9�N���Ci��7`�f�Gۜ�K(yyA�Z�ت��`v���GȔ�s� L4��i h���"������$PI��q]v-ܣ�I!B_ݤ�Q[O�Ĉ˅�a5Ԫ�Q9�C���'UH��i�(ԅ0@�8��)��R�	b,���T!)�î.$���=,8P��X�k��s�\d3'����z�L��.x��',�`2^��e�Z2�R5�j�0�ar�4b��T(��9�p���Ƈ:�t�z���7�d�m�R��ɛ�`���Eq����׷2G=�q�����a,��*W��%:��1l�D$�Ɂ{�aq�'D8>E�Q����E��4�1E��^��l%=���?��m�d(��~�aq;I��.�=�b2�N�W��J澰c@	�9�����ڲ0;���H��-%>DIq���O�r2��L��{1L}o��*�t��,?��n��,Y�VͳCE���V�8(?Kc<t�h���,ID0*b"�'�юq�R�˿3�kl����f&�R��>	o��'��-�Ai�s�TArG����c�F�7���� �9	�[�҇)3�,�2mi(�xL:(�<�T�K>��Q!~���,b�.'��݇@��{'��X��
ǡ��L�1A�?�"�gR��w%i4�v%�)���/� ��a���&K&┅9��z�p�<>� ?ѷ��xf��\���J�^�R���Q�BBla3ǀ׾Ee�?^hEx��Q�*}���Ī�����V��p�P�a���?������f��$��E�����Ʋܪ,obUY�ms���}(�ZU���3�&�모䱞^��1�7d�WbY��,v�u��/�#e���(�/}rI߾F�����=�pp�wU��]>�gB�{
�U���e9����bmc�Ϛ[�4���U�6�AXAv�<I�E�aiq>1���T���{��yYB��:��FRߋ1�����T򻌉�bX9K�W��o ػo�Vqz�;��m�������1���d��>�Yć�K%�9iS��$Z�\���N�M�R��{���m�������ҿ�x��<�sBI�'�=㝛O��5-}S�	��10W��>[����ۏz��5M��E�W��pFe�[���4�������ÞyW�u�~ut������Ko}x1��`A]����uϮ���+���k>uUI߻����=���e"��\?o��{]�;��[�7����޹⺻���ɕ=�wI��ԴʚI�+4"Rw��Es�u�S�I�3������^Iض�q��������<���J<��������
x���K,@0.�0��������G�E��m1j��b=l�S#����� ~������B8n�Ut�[G�`��닑d��g�+�2\���>kq[x�?I�)�/_2g������^lY�|8�P���6�W����ݰe4�|�b	��mu��Ⲱ(H�Z{���c6G�~�`�U�����ἼC����X����~��q�kzKN���YKHc4L��w,z�S��P�o��+����ߌTe���a��8��R$⼪>L���1.D�l
}��ltKf�1Nf��Q+�n'����@6����J�}�#v�1�_�I��9xӊ<�$���y^{"����A9?���W��g�p�lLFޖჾj��5���Z0<4��j|�&Ǘ�Nl��	X�HH	}�:f|NI^v�Jg���g�B_�7��bIV��hOU�5�?I�h<_�;VU�f�Ú�
kI��ZZ�ٰ�ޕS98���̅�F�=\[�$ba�9әa�����}N�>�-�
cwTa�E���G�zC	Bp�t�%���VofJ"۪���fL5���R���
+A�j�"�)S\.r�;��v
����CA�Z,��le�H ����h�!W� �\�7˿J�Ϳ�!���~G��^�S&)�e<��V�+ĩ�#���~���WY�P���`FKK��XTgw�E�8�8Ü�2-�영����e�xX��>���P\$1���a�)�� �,VNR�iru��8�)?���s
"�HɂhMg#)?A�-K����M�&'�&@a�*���G]�����d1(	0�$��$��RԼ�ͤ��_�o���� ƨLH�=M7I��r�,_0�m( �k�5ާ�M&#7K�BN��R�zu�t�F��#���h�*e3��fp��bz�	&Ip��M7��9�}S�8�6*���ň�S�D)�-Ͱ�l�bҁp\r�,�%��E�3;ۆ`S�n���̘��crbR�L�8�PM|� �
?���i��l̥��C������t<^�Ya M���b��GNN����g�I�KO���;<(�Z��j���8rD<4����?�	ZW�x�X+g����¼������.؍H�OF��X�8V3������!�]��ɹ0�%&��5����cf��N�ˀ�g�53n%i�����Dx��āC!@���y�������Nc׸A,���^3�T�����Q��ݙ��4<�][C�T�
vG��:�z�|MJ�'�0::B��ž���!� �#��:�l���.�Kp�y�"����CEy9L�����8�2I��"*[ո͹z#t�]n/&&&��+ ͌��o ��v�d�::{`�ڡ�r������HнNj�����1�ν�^��PK0��'������Ѣ������)�Jn����� ����Q�;H������^6m��b�u� ��Y���pn����T�``���A,OM˥3���s����z�58f�r!}�X�E�`� �-��%�f"F�V����ŭ��z� ���py��P(�,��WA�]���<�x��G�M�0t8��Q�z���(/�$�"s�*�%M��+��6�Y�u5�J>�Qbő�Dؕ���`c�Ew��^����ed�K��r"����Uޒ�)a���;��`m~��9�9�D�+!����'!~J�Z6u�fT�ƨ�L�c�֡(j�U��|��6u�s0�6!�;�M���#Ӈ�e��$�iCU�^l��� ��B��i��������� �������8>���I/&�F	!
h0b�1��#%�2X�}���_�:�7����@��B�����H,�,�[v�q��D�	��7�����6��.*�$�3��Vs�s?��K��QBŉ�~�!TC��8$`X������:�M")�������>L#	r�Bdyr�@z��1���xz�`��]&Nm+���4��SQ�M��Z5��qZ�ʪ�WW�|�0;}x���:�g��a��
���k_*I�����Ș�    IEND�B`�PK   ���XhT���� ċ /   images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.png�|y\����Td�D�+!*ZD˴qk�J*E�B(�F��-��"d�V�j�s�!5hE�(��}�]gD��<�>�_�^��m���s��z_��u�3~�5�7od߈�`6��(��`60ƪ���/�싿��8����������7ت�s�`v�F��)�����vCQ�������/a��Z[:�_��$dcoE�a�`x0�
�u��}�R�8��w��`��&���`>�kq���x�i����-�S���q�A�rg1#u�]�u�\��ʖqѽ��D���A��뗬M�N�Wj��S�1N�0�����^a0-ⷥ�^2�;R���@�z����f����n��=S�u��x^����:v�5��+�5����;����w������;����w������< �M����R�̼��CwR_y��ح�|2��t���S���]o�[��}��C&-�Y�5�	Y|�F/	}<W�|i^u��b�ud�MK�e��W1�F�]����F�I�G������&Zꅽ��c������7����Ϳo�}����������lY���и�vKr������?���dfE-���aƪǛX�nd��z��"��&�99����]�ʎ>��4��u�8�O �d�%���	g�}��&U���x]a��{+�;;�٧xՏ������ZB�����A�ca投�B��䠏����d�������l�i
^�QHȤ�����[W����9�9�nj賍q����#I�_��Y�6l���xrR��Ӯݙ���\�/_�Ħ�:�|lB¾���FB�q%%r��~ۄ5�*����i;�)B���q`�~�*���;gF��:+�l<�'�%o�9�I�?�w$�+j)��˫�,ѺU;�_�vRU8������Z̕�~�!rMG bf(��ْen7�����^ &F��}��l���^
�ŚU����M����{���M�yWVRPPP2�9A-�s�[���4<��ʕ[����!ܚ�v�������lb��ˊ������x��e���fii�����C�{����ޘ�׷�u}xv�n��Z�iĔS���߄{ƣ��yL�Q�'L�9���\-q|���M�99G'�~�)��璛����Y6%-y�c0+� 6&C��uO��\v�zK�W��a���[k�L_���g����sRv��Ǒ<St�fF��d[h�J�l߯}Jv�OP^+5+KԺh�J�`{�����ʬh�}{��٤]&��oү[gnjʣ#�w�f(A�N��ŕe��>298##\Q�jtS}���$Q���7�|���	N�f���k�:9===���h<��uA"������o�aDј��\Y�v�
�U]�*�SSSsbb�≔C�An�U���vRڑ��k^�7ݺ�3���k:�H�WllB�ڔ�>8xnۏ?�{W���o߯Q1?\�=\<m�6���˽������^ϫݧf�^�L��@vp�4��p1���5�u%�m�B���뿼��/-�K۽����I1��$�]��WX�֐�J@���Z�;hTp+-�M\կ��r��Ü������~]�!I��0?��f���󱣃;��ACC,��������l��Us}ͳ	Q�J��`�mk�������\gF!�?77��au��[�I���%6��76oN�.?��֢e������b-��3��&'�sJ��{��p��;v�����R!ս����r�#̓㐣sRY!«
Φd����hur�����|r1�;�l���M�Qd:*��D"���rdY6g �&���^C6dQԪ�U0�h�i/�^
��]Anb�.��������?y�ĉ��Ϧ��Q��[��;^��\�Ӟ�,��_;:ǉ�w���>>"!Q�.B�+ڕ엘�H=қ�w6�t�,/X�	�}s����6Zǌw�ڔ/,--=OM�c���-����A���I�'z֐x�;�\&�KܜQ@R�.FL�Fʝ'�͇ۋ����b:R��Mi�;��)��L�� k���;'�MB��m������[@~�	FٽV�S1��Y��,�3���-	�'��j�Gf��ή��Q����RT`	l	�^�4�$i�]e@j/��~^��QQ�)�vLJFFF|I��.y~W�Ǹ��{�e��i�������335�M$J���6:]�,�4YZ�H���¿�n�E��SR���eV����T.f�}v�0�ݺ:C6��G!�Ĵn��p���Q%���uuuN��������/�Mca5�=}��o�G��~+!d7$��#��H��n��F(W��8l�d��G�V�8���.���˺֘�4����ݺZk:������Հ�q!r�,�"0����l����D����|�9MG�A_i���Q3Z�ɄP��������y=���7��[����㲑� ����Ӆ���c����m�/]�v��{�.��hW!H�g������O��:�8C�jr[a�XwM���=Z��;�vG�ef
���h�! F��-�a�� ���d5��0�!�sww�Y��ʺZ�x ��T�|-��KJJ[j/�.��h#��N8��JTfm�y�?��s�OԌ�%x6�Q�jn�'.[�TI�	�]o������ͩ'x/rߏA�-��6O�=�&�z�x��8_p����C;�ߣ��E�/���Us9V�ºH�o'��ЭoM}C��2�
m1Qd�c�b }��~�ª �	��'���-+>�����d#C[�j5)b�ޅ���e���G���V�E����mQ���7l狧v
��g�v?2b/�Ĺ�G&k�l�ׯݔ��dIOv(2!��jf����
�Ľ��h G_J��?��@ �h�Y�?�m��I�^[�{`|]�I1�ʻ��1�N^^Z���|���@E%%Y��j�^}��`q�����J �@��]8���fn�;N�'����������v��ф���1�@pnR"�6���O����z�Z	��<f��8���=�x#/���?~Fޑ�����8���f]�۠����SQ�v
s:��%E�%���tF�.\:���I��/�Ja���;[=r$ܥ��n[���n3ʱj�/�hhnN���Ɯ����oC!*~��A.��LG�[	h子2�����Q�uj1@F�!C�=���|�ܻ�.��5Y��\Z�c%�@o�:<\���	kD�<�/��ikk}'���o�!�v��% !��@)t@L`C���\��L�V~�X<�;�
V-�z�Ȇ[C.�?��4�Q��o4�p���-�Y�	6�cC3�V��M��� E��{ ��P���-¿��=�6�"�M4d-t�L,���jB��R����D�����Y�(	������$yp��+3=�<;�Oe����8�v�����Y��Gk7�!7�m�w��i6��D퀁/@�!��K�[�mpHyP��E�i��B����E�#�Kz'�nr��>���W7�?�]� >�������˓���F�f�LZڃRG��<W�~j���
2���]&�I\��^����E�x�g_L<�O����kF���k�a��?�4�z�y[��&�?��9ui��p�%'����uA;:Zͭ)K��Ϸ��C���X���NX>�P�D�:�bt�����#�~Jv�%�4�S �� �.r��^��B*��S?��!V&�|����(����2�b���kq��%�s����^q���T*?#jjj
t��O,�fVL3)�����F#��#�)�Q �Iѡ;��#a1{a�%b����J�|��q'���>���H	���Z�!R-[)_ʡG�e�����[�kܧ�X �թ-ɺ2�V��`������'e��i���=��c��f(��E(�W��sW=IZ��!x��g3�|��}^X(A϶�q����Uabj�*�(����4P��w������~Ϟ=kpeWt�?2ӭԮ��{��E��Ln�e��uD죭�(����KT�3����^:S)l�99)� �A�-�{��Π��?�í�կ��?~���Η=���CP��_�����"kFA|(��˿����dXN���m@��|j&��ʦt�8v�����r���&�?�OZ���lqn2�"��qf��r��n��v9��r�{F����wC��� F?*s'DN�z���H��_�����2L ��-RE�D ��m�	��8Pg�� �S�-�4�M�_�۾�
�7P�?V�p`rrr����"B�K��e� ��T�eg*#����l)�YR ƾ-h���U��c��xO�����uR	�8�|�KlT*�\�Fi�A,#U��@|"%&n�rυ�j�.�Ifs���qB�6��X��vC��#�X�n޼y��M�
���7W>���[%�l``@͘=fɣ�ň
Z��IW�l=A?v=0�V��?S�ɉ�
J��|TR'y��U4�jSG�JgV��ԹM�ʊ��/_��2����pE���p˳�ޮZ̈���{��1)գ��գR��FR[��r@F>I=�M�_�:ܧ���S���CC�ww��dX��WZ�Q�8�=C$\�� H9R�S�I�^i��U荌����39��s���`�d�Y]L..�����I���M9lkR�d�������(...`��)�CW��m�����{�߽��Χ�H�N�sǧ�N�0�);�:��^��V�WD�c��������!AduP����zR
Q����a���[y�z��sܫ�A�ժ�0(�I5?)�[��b�eA�X�#��G3-
>�����p&�rJ�o����%ub�$,��Uy9�=���c��׍ǚo�R���]�r�ލ��e��Ӎӭ�0^�/�+�,_7s��e���+X���NzN({2www'��5>e%X~4�d�ڵk���C���G�B�t�������r��囵tu#���x:5##��&2�nF�΃$�n�����R�	��;�ϯ�͢_([4�=�)uGT�D�5<��Y��2���=d�|��2�:�}�Qءgx۵�~�̽��h���ԟ��H�K�����⤻IZB�8y���PEP�c4 Y�N�g���i�j88�E]��9�r�I�]��e�Ϊ撩�Y������婎��ojj��ۘ�lIK�Dw�w���9�&T�,��))0��v�z�j�}͡?W!=\$���57�ܺ<�,��z����	���� �����Xj�F�F��_-����h#���'X�s�,�E֋�-��I?�#  (��Ǔ,�q�9^�֔��/$R��4� ��?6>�*=[�8��&hib�Gxx:��O���M�/�zӭU1��ꇧձ���7d����|�� �`0ã���|ڹl3�֌T����sM���#�&Ï�HK�����T�>���Jܺtqj�آ��G^Jj**��[o�z��y໧�؜r�E���x�!�������\*�XGF����u�A����6QS<�#�w�S}[H�/��YlBn̤�^2$S���B��C)��1I�d*�f-"��ɕ*�nn�<d�S;I�G�W��?��C���z׉�2٨Zl1UϏ�y�˖���HJdu��1�~�rJJ������e0}ю�j�s-�v憾��ٚ�0=���iC5�c��s�bލD��"R^Ϻ{�l�a�S�e��ZFFm�yTO~sdnU0�������0/�����}���v]ASs�y+
�<ON�O��n��0�l�}�Νb�Z9B��x�����H�#�g����S2��5�Ɋ��v?r��*��6�5��7�]m�率�(R
���I��^�"��L����##Y$ڝ�mLVOS0^4Wj-��n�M6*8���k$�7�<5Wz�D*[/�q�n�2�87Ox��S�i2�3�"DFFVs��	���N����d�#y�����kը4�H�f抗�j�f������v��z�M�T�aU8�i����2.:j�*�Q�q�}���r�s������Ʈ�m�����3�v���3�]qBT�,���u�������we�_,3��r��ܦ�ӭ�R�Q�sb\�9"���y���Hj0��jL�3�pv&�\��*aݚ`L�%^�M��Ή:�}p!�cl�K?�K��z���s��݊�á����J����P}��{0���ȸ�UR�ŷ�o���p5���T�?xP������s�[ �	2��u�̦zXdm�e]n����S{� x?�Qov!��2�|QؒD��"����A,
�I�cJvuR?@P^�o�娭0?�(.���������Q�˟�7�
O�QM�A�Ņ0���  rST�:�<̿�8����:��CWW�e��ݟ��+�;�N�ZGRx��E!I���f1�����8��Dq"!����[~�U�$lb'�@�G����d�E�����6R������pȆ�|n=]BWH%�T�3�i������c�+_~�B6z�T�Unn��p����!2B���7m"z<�����s����!������{8��B����qo�06����ʹ_3:������'r�Xt���39��������*���,����o8:�؟8~�833��ww+���1oxsO�03��(�K�����'����E�s�.�aY�DJ���0v���q���R�Xk:���E��
����Z�0���>��uuu!O�x���C�^~����CA�]��@0�c�Ν;�&���{<�<D�@�7g�̰�9b�ޠ��q����!��͂����Ό�����h���w�bcy�N=���4�y0h�|�8a/�&�]a�:g�N�g�Йhkk��r�좙�,������i�����A�a|��a�����5�[g~?�OmvCfLsYqA�;s���G>;q�����]߇g��DB"���%���k+t����(]�t�T���Ј��xUp�m�\�E�g�'6������.��/�X==�Wyyʎ�ӟ{ݿ���d;� )���l-f�>+�����7����&1��l����x䞟g'�$2��0*��߆ey./��zz��%:�EǸپ�������,-���{aK�"M<f?��Q>��+IL����\�_SIM��s��21I3&���	�5�k0�]�}��Μ��l�UU	�g����($QV�V���rc�D���e"� ���C~ʒ��9�����)�&9En㘟��>?U	����8�:Ɇ}��Ri��Rdew��.�ˈU��n��e`����R�0_	����x"ɴ?�|��W/�����D���?��������uH�x3�\�qDD�����d ��$��pH�Kٍ^����ۇK歁1I��ޯ�v],K�}��+W|��� ��4���R����"��=��T�/�c��JKw�,u�tR��x�= lX����:�S���qpp@���o���!������C������B��0>u���OK�`����g����CȻo[{l6646Vf��{H��<�����{xc�	gE�K`u�_z�B�i���� �:!�Q����W`�3�ی���K	�pهG��A�K����yB��dŞǸ�?׊CA8��:��y�����If�ux-==0��X?�Ą�}��c�g��j9���K����(���"��Pd �J�7ݺ�-_:ܧ� ����i��J�����1���QA�)��֛}yuUԼ*�yZ��u����I[D���=d<M`�Qu�c[�w�;85�q�d�{���YH:Y�c)���y�� �m��D�:�aT\��U�vr�%%�ggg�}�l�����L[_�˗��)$EԄn�gI3sUm#�]���,�H�H��,]�Ƣv�d�A���	�b<
5��.����a�v_�kQM���H�ud����,�Ůĥk���B�� cCCN4����CYכ��J�Q���eܨA��K����Z�UZ�|�tqq1�(qGN��c!�p��˾��E産C��* ������C��������<OM�X��rnG�M{��--QMM����

(�!���i����Ec���5z�4J~rʹ�͒:|$�{㓔���N�с#xo\z�!�6�
T��9�5���0��7nެ)�+�N�%o����EJ���XOm����]<��QP.��^9���խe��5ݱ%%r�܊�u�����:�RN��'��2p���+KaBa)�%�\�����p봸�=�B�� �����cW�C�Ҝ�e��l�P��"i�o?�������/I�����,��T�<".�X�p�һp���*U'�Դ�ۉ�B���כ�oF��	%]�H`>~���F��k�ޥK���^�I�̴���Q�%e�uأ�*J],��2�����~u��q�Z�_#��X�Yu�Ȣ@R�}��C�/@�qF�:Ec�k�׈|G=I����G�Xl�y�:2:wZ�Y�*�Cð9�PL�٨g���"��|��B�!�Y1��u2vB����lVgz^�?�'X�9HX,:nϏ�Rvo�tyz9��u:zqF]&w,���|"�uzz:��ӷ;,�3/ف�4
aꋥ��X7���"/��?�`��� �mY��I�F�ʻ�ө�%XHgz1��3C<�z=�������M�/n[#��%�$"n��j�kew^�������X�#��v��8��V��WM�=J:_s���ANV�;��y���>-/.��h�B'�)�� p�t�7գn�UsK����)6LLlv�*��̘M��&;��]��		␨�
�0��aW�.Q�Y�'�6Qc%�L1R�V�ER�6��������CB�d��|с�=C&gg��z�y�������I�A;H�(���r
O�y��	�0l�u�R��:��P+P��_-~�����"ؙ���|�׾mmmZ999Z�f rv��͞�/�a��uV���)@4���.]\@�9����q���]ee7He�3�l��
�uR��������0d�h�����_��}�Ơ~-c�����7n܈����>w�-U/3x��Y��8�h��:.�#~^�ok��ez�L	.��+�7�@��E�ĹI�h+2=���tq�!����+���#��0��]J�?�vHFN�d`ˈ(��T?�4�Ƅ�ֲc�5݈-�d�3�e�"j��J5dv:���$g�"�k���X�p5�,�Z��X�:��!;��͌ҥ9h!x{ZA�C��ސ�ɫ��=hX���%j�	斏Ʈ󉘛���s,َ҉�K㨬�J��F&` �o�s	��Zbe;Y_"d���@�b�Q��0��:Z����An6
2t=O�?JC��I1�Vw+�pJn�l�BMZ���v
�M����$ J7Wo���_���O�>m#�Nʀ��	�M]`M���|��nSDqy����%J5E�2���>��@��Ȣ�=�*�]����_� ��^ֶXq�W$���n��⼁�6���ظE-�Pԉԙ��:`���[YŕBvq����i�<�6:1q�yd��h5�/�Y�<.��Њk6B3n���Y�܌��4 #�:P�hԺ��Mi�L���<�q���[�W��ᦦ��K�e5b;����~�'ʦ
�5�<8���=�AR����P���T��ػ�xzQ�o�֬d��)oɳ1�׸�;�jD��

��أcccr]�0���);˼鸹��� K?E�Lx�9�=��Y�bH��4Bg@�Y}~�����B"��ZO����w�ޤ���j {"k4n]H �Ine�,;	�� B�{ooRm���uxHˍqYwV��`�%3_��гx��FXP?�ۛ�+�%�q����e�Da��z�~t/��L���5�3��>�wtǎLL�[Z7m�LZu�1�k�5,������wd�������)bB���Q�$�~��%����LiN@���^!v@��-��ء�84�;w ��>�F�������Ɣ
:�������/�Ə��r�V2#�H�5H��m������ˋZ��[��x+��g��>e�v$=�8Ib<!�-&&-�:���у^ޖ���G�/Z�63%��R̓�!Z�k��P"{�ñ�4�i�g�S����M5�jt+@�7蜭
9���D�.y���A��ao!�L��|�F.s�D���F�!ȓ�N0VfzL�J:�����B�l`�]w�p�}S�����4�KD�����3ޯ�9F>�A�鐺�ΟgG D������Hۖ��"�qi{����܍�!��jnOv�Yt�?�)w���|"�kvv69le���������q��v ����C ���}�D��0!�v�x"� L�����cb��Y�/�yu�㶈x!>Li�y��%RY�Wx��h�'
�;��Jĥ�
�}���:�Aڣ�`faIҠ�95�2�n�4��ЗH����B��WWø_z����iS4�ĉ�q�r���u�+D��s��c�A����h�KK5<�D�^�=��z�OK�}�UIVbGC�	��r0*3�b�QY�wɲsHX�����TV�Qؕ�Sͣ��U!�]����Ͷ��~?�v���� n����d�P�̑n�g#j����2�d`SI�(��f��o�*�ink�B�r2��܂۶����,&n�M�,��Oǰ���k=���'�gGa蟀�.�vUT��&��X&u��y
<y�%yR��T����VN�}����P�1�1k%�|��46�ST�:V/��ǔA�A$j����2�QZ�&ɁFl��¾f��#�)u��i��K�;�Az6��:�*3�7�<�;�`;3���Y�s���uA(�v	��4�=8�ʾ��>Dn�
j�E)`�|���!Sh8��X����hD���
p�����g6 g�����J�(�k,֑�{�&���e#�HQ���u�� ̻0 �E*1��1��Sh}�wt 5S���q��t��]�J���cSRP��WŸ����	f�:��G�4���_鲐�?j�꓏��L��Gb�uO�\���r�M�)ӄ;D~�	5N��A:�����M��yT��ma�sLj��&�zz���Q��6G� 	4����MN;`"~ZqJ	+<^�r��x�����/���9�pw�qP��{����сO~�AjMMMX�\YSSs���ԗ{����)w*@
Tz��ڰr�R&�K֔�ԑ��fj�DĶ��3J��p��'"��l�q�`�P�|��G�^�H�d�б����ZU{������~&�J��2#���6����S	{'d���?�mi-�#��K���'V�>H23�ۨ����a��l7��DDDh�=����b�Ce1�}��0���^)�G�<fPhݼI�h6rL�Ja��xuW��.��Y"j ��x��2�6J���>)�gQ�V����r�w~�T>צ#����#i�D~���¼���x���w�O�Q�d�Mu{�+���,W�r*H>�� 3��c����
�XY���� �{
X��=�����f`���E� �@�.��$�5�]�TUo����FY��o���Q~�va,��&��<+K5G�rf�vr�{E�� Z���=n-���RSfT��g��!��j�	ʚ~�l
W�a(^ڱ
u١z� ���' �6œgQ���y+`k` ;�F_���񩪪�<��"%kc����Q
�)dط��χ�n�`ع��.��Q�8�8ر�hW���@����
�e_v�
�?�L5�vG��kg��p<b�O�W��5OhSxx�o�F��V�\���<=]Ok�
�k6�S���yFF0%˰Ə��B�^\>dH�=>�j:�q���.�	�̽�>�*�PB��ѫ�L��x��k&�L��O������Φ8�����w�i��<`�8�pSF���/y���Ѩ�J����J:�]<���,���x��×�1n�ŭZ�������A6E<Q2�j��u�O��h��J6�z݋���ݫ(�zO�/�/44�R0�����~=pP�hkadHU�`�Al��Q�*�}  5�+?~\GWm��JFb��BC�Y�.���MX���H9P
����<�XEy7n�hV��Ի��ⅈ���PH����%�S_Q��TJO���u��c�GG���2?(�ߐ�bE��-v�{B/ 2�L��'�]F�`D Ea��2S��pT�Ӕ�����X�3�J�c�~�@�0>E� �P�?<\���������I[J[ZX;��:��DT���C��@@S�%��9�`۲��Rۦ[4V
�	`p�H�VN�<ʘ��{'��c���^�խ���GU_�{::6\��H�L|]4}:������G^�.�8+7��r#�1�݉���ʼ<�D��^^�޻uF�{K�X�	/�L�?�ޏH$�IqE@n�G��!���M��	����&�o�ܼO����u���_�%��q�������$��x�Ow�����W����W�&j�VN@��WX�踞����U�c�8�>0���@�w�ct������7��9�\D��r~o4+$��kAlv�/.D	�E2�hyxx��O-����Yv�T266FZ�1�V@�9�3����&��J��L����IO��5ݔbP����7�����=��8n��-��̓���Pj��l@�Z(��쪁�ch�V������\�h���իW�5Rvya|�8��s�6� �r�Yݒeny�By E��>���V$G�]6�S6]�˽˜ঈp��21}�j�@.�N��Ać����ς���AG�a|�'�ƨ| �>�J~S.)��%��6U��ڿ���OQ�r��Uកg�cD���GI�C8P��P�/Û�/E��s�{�h��c�!v��v�#�N�b�@�no�֜@��9v�9�퓀��� )G5�3�ފ �Da��_���9swf�t�R>�'�)�R*�6���sb����

����&@Q ��8���Vn�X��(K��]@5���mG�g�q���b�{{�o��d��.���uG�ЅW��U��ܞ�,�Lj�B���Z�ῐ�?G'�ھ�\������K�X�k�`���8\%Z;�C�䂚�>�4ee����>�9�X0&$$��=cg����߁�{������î�9��2�{���k� �)W��mu���z)))�0�e0�@�����.��b�e��H��b�d*'Sѣ�O�Ao���	���򳪨���AU�njlA�˛�e\B��_R$0G�k�˱I2�ߡ��+66���VA`y�⎺��.�ꜳ��4�ѥ$t��.n�ߣ�c���:�N�����A���E+� ��S�n�r�b4����K~�3=���/�aFU�ъ��r��-���Ы���n�1�}�|�5���"��Kl>�a#�YhnnyIm |����*t�1E�'�r�x��ȆXH�����B��:thT�sB�w���K�_����
��BB��@���kx�.��R��U�:�mܺ8Љ5d˹���FFF��Þ?��7�.F�����(�FA��ϔS�v��E���U���@G0ԯ� �> ы
��7���6̼��t�ċ��g[��:��k��:Ŷ�J�Y��}���c���'��A��{��7����X	���`0��l�T�%F�P�̼�+1��r��,�T	��-,,�����A�:�42 ��뼎?��9����D��FQnq>�f%���*U�"��|��^��Hq��Rί��ji1�:������L�H�Ofz��<QX��Zzzz�ʅ�y����M���?%��m� ���x46fO�H�\�~ݰ��W/ �(�4Y�4�F?Iыq_����1R���葘E8";c�04�>�+��b��s6ғmvvivew��b�0�ʓw��#���~y	�{86�����u<	>��m����7���}jh�7�l�A�e�V)�#�}�Qt�k�&v�=8�SD04�vw5�.�ܖ�;BJjJo���)'�`����!%�ݽ���=�-��9(���!yd��X�mص#�t&����A�������#�fdϛ�麻���3�S�x�Q���/�H�dmS��wWh+ڦW��]�G6EGI�帖���	啃dr���<2Y����x�	:GV> èV�N��O�H�.3 <ѹ���Tp�'ORΙ72��+sEEE3z��~9�{<��|�$�*UYY��-�t��v�Ζ;��={v�g+qT�L*{�P_��y�a����.�O��	����vS.T��]:�A,�F�NR��qv����xI����r��1���(�u��;�v,�Dw.�����R�b����u����F�G�tK�T�~ѣծ�(��EҖ�����T�/}@Q$��m��eSZ���[� ��3H��H"�4+��.Q��7��
���@����PzKQ���1~aa	ۻ�#���ZN�m5�!��"�G;�
��tZ��_�Գ���w'̍� X/�.N�#�~/a`�N����εs~,�pٍ����j��Cg�讽����\�h�M�A��x'�1\@���	�᪞����Ћ˒���9���&Ƃ~BGP+WFD� :����o� h!R�{�-�#@� F�Q��;�y�P�Z�����D�|�AO�O׊SB��(����h<@}��8nE`li�s~�&3`�_//N+�R��m@���*��U�X�6b%�t:�%5袞��(� �#����r�Z����Zq�P��?�\2}��f9���.��_	���� ըe+����aJ� �|萐xc������G`�T`���0
��T�^�F��������o/�ɀv.G�G�d��?{I�V����ۇ+~��5$�P�<�H^����;v��>`f=��y_y��=B�� `������/z�:���9�Ά]��Մ��Jщ2���gm�	L����pr$����+��%(F�,6����Fm��@�mQ��gՌ�5�/���rFyN$���#@����]j&sg(L��%�&����Ǧ���u�?QeeT��1X���X:�Z�o�������Wj�i�{�Y�~���F[�AZ/����A�:y���C�����Qy�H�cS��y�."��}}}*����$D�������s#<��EZ�����sM�.);��:�D���υ���7I/we��w����G�~�U�c6��~<��z����6��ƛ��C�~Dg���4v�Q[{_�?�o|4�{�y��硭���S=�Mt������M8�Ǎ��$�bZ����Bx]�#��~�ć����D�v;;,�@E�;�x���{"�o3���'c|��i6��&�z��<ʽ���1D|���v�m~}���x��4mL+/�-��k�>f)B�|�� p�E�W�kʼ.?K����$�U-w�����b{'DnNE��Ћ:,�Ѧ��e�Ś҅ {�t�3 *yDA�Mt,/v����Р�ݤ�A�:��������4��*�/��K��%�i�2��өO��a�F�|9���J�Erl:�ҍ��`���:v��A�K?}�">�%����*��!�O1Nk�#�z��{��$3���[�][ڑ�O�A�loLs8�v��L�D0�4$�h@�4��9jO> �]m�����R �#-��E�Ν;MR���ӂ��0�@1����f=�]y4#�X	t�ϳ����������N)(����wov��=qx9�/��z��z��Lt���Pey:�+A1`����s�Nx<Y C�;��[`f�1�z�oo�3���[�n.]�Z�_2O���vb�K
�c���=77��z��_�}�?�؎���������7)������dքH�kld�ϵ�l��!m���Dz
lW7(8�|�1��dV
��޾ͪ{�1*B�288X�UN��X�Ɣ��'�;��Y��_i�ndccs��l1ǽ�o��.O�}������b��6��dv5[f'��2�ij6�2N��=Ϟg_�s���\�	~=�����Uv�ų=QX�@8�䙇r���ɲ�ȹ�?����SH���`fjqqvm�ŋ�5��;�|���v-??�e����� s�˗�X&i"[�]%L�o�Wx�}�I��f�~�z¥/i��p�I���/*xΔs�1�Ӓ�h�lIe4׿�z�-o*�������#���XmC�O�.RU5N���cץ4�Ь��V�Y0�Ž���n�x|zZ��A������w��}���1K���$�o��6E�>��Yv�R=}ݑ&g���q�o���F���4"�Y���N���;�g�����t�u�>ncF�ǲ���Mh_�d���Zi�N�cRJ�6����r~����hwUa�89R3KR�^��5biɣ�9;G��] �@d�B���Ǘ𷈤+<��		��z��uz���Tp@Ȳ��^$�_p�M�q�����+7��k ��q�^DH���"�W�KZ\\<���U}qq��?�h"�b`qM��`zZ��E�_��20�@�ƺ-�/�l&&n,�T�����j�AG~u��器�y*�s���z;]̰�w���XŹ$Ϲ�ꏏ�Ů3�R_K�Ù����O&���rȮF�ib��bbڈd���ߒ�T��0� A����0�q�ܚS4� 4ū�M�:Q~l֭I
� �4ИFdgA��$rt�G�BGC<u.�ᇆ��v¸p����]�9�H�8����X�5��	���8d��[��~�M�W ۀ�����&6�RFaa��/��7��/H��T��񦦦^M�8�M�~Ih�J�d����g�ݡ�Hh���a��{id��~�̅ό=f/��c��u�v��,�2���O㴍αL�%n�E�a�m���H�� ��{�f'����L1��I�s.���|� ��F��}dL���kW�f�ad���Y��q���a�4��=F7�?�d�dD����)A7;vip��1�Gn�DwTB����x
���j��2զ!�tI΍�,��&2�i�,�D���v�Y�ﱕ� �O�m��`[��ۅ�Y��YJ�=�\Br�*0�<p�|������iڶw	��z �%pΗq�mhh�K�K��Y�	@Jj zL�]�t	�a���		��tth1s���!'MLb	�,g�TPp�(7���Q
.B�LG3�u�oJ;g[@��DY��=ʯ��o2��	]n���S}=�j�;��e+%i��Ra�w��v���F����J��C��!���l�!j���:�O,�2�������۷��-����I��)�v�~�)��1��w�d2�����V/���8$Z�̛�2��x��֕I>:|��ev6��M��D���9::�&�c��I[X�8�Q���){��T�cWY�ʮ^b����� �ޕ����I1M����o�U%���y{��� �y�<~�Kέ[~���ӷ����@2�yp����7LT.����_D*�D��g.���~�g����1S<���)[���0}�����e�m�[���P��8~�̀.I����#22VT���	���132�6Gv,M}����*�㘽~�}VZ:]�+CEL0�H�qƽ��T�S�y�i!��|Ȥ��*�v�â~�d�ê�<{�ۣ�v����{�fY�@�eѭ�[d�u�s�1�,�\���ڎR�[����|��K~��xmmm����ׯ�2*�	����L���{	�a��5i�1����i���*��m��~�E��o���?iz�m�}(Z�]���CZ*#]e/���I��G2� v�DS^I�2�{�n��ӧ�B@�R�����9u
�=�Y�1ʦ�^��IH��D������Z����x�@�]iLѥZ�ʅ(	��o�w����4���^�{�QUS�>~�G�e0�V��5U,���6�i@��[�ݧvĢ�s��UP@���.h���տ��p+��!��	w�ڵ��a�%�ג@�#�d�t����2��2}?~���ƀ���`~Y�i-�)�7@�&��Wo�VE�[��J��6t@�����yрf��e~7x��5<M<��=h�{��ly+���t��� =��mbB��6��(��~&�g��
�.�=>��m��}l�s�Ƥem׿��"��pJ>ML�dp������Qq�%�����@��l�/�۰xy�v*��ZXh@!�w:;�����8����1����f�{IK�hJ��˄����z���'A�׼���OHH~�ܪ�ȷ��e�G^�d0n�Fd��.��7��l��عs I~1���ð
��{Eh�@F UW�Ux��4NG��A(��[M�X�Ƀ̄����Y^��-�J%A�U�jy��t���x�c��`��,��bbaa Ȥ-����|�P>Y�r�wö-ws �r1��3��z3��у&%�����������k8)H��Ѯ�q]�K�0�ͳ�9@�x����`��V�@����QU]@P0��+ `!���}���?��4Uo?P5���b��Y`�ɘЯ��H⹊�\�^�*��x.!!a�J���&���
�A����EkUqpȖ[�1���/z�1�"�b��?����a� �����{6��*�����}��s�U�h(��0F�p�V�\u{u��o���ÿ]�_�����?M����2,M�ѵ_�_Q��jaٜ����(0�9>�q~��zLI��_1L`DoJV�G*�T5��%��F(�'Ҝ�&���Ǯ闸�g�&��'�I"���_��6t�c��q��*?Y��+�Y{ěVYhY��q�s�˰��ΝsY�퍸��6�[o%J�HJ>oLՃt�
�G$�l��3��/$B��%���dΓ315�ĸ�7<�t��Oi1X��Y>$���V4���2�)�UG��I��ЍQO^�� AW~��.+�e��a�n@���/.��B�`�QWW����؀fF�Rwlp�x���j���d�
Y���,�b���l�C��끙'�g�<���3O������qtI��6+���~�p�Sa���{�8l��r���u2gv�����������-Tɚ�*�7ک8� �}�Qf<vd=H�4���T�#7�#� �+]�a��v�ݻwG��d؛���$ &VP"���4��*M�R�����87	_��X'Z�}�į�l���1�O��t,@��x��n�s�Nѹ@��z�h���>��$R��jH�;}�=�Nd<dy&dŉN�l�]�	�hT�.:G��a�Kc���a�g���Z��M��g�StS��Q=�w��irLW@@��M�������D3Z!;�J�Yy�U+AV���I��s������g��	��m*�A�]�e�s���X������Ů�����֛�S�>���;�ž�J�TDYCZP�d	�-�ز�Ѧ��&Y����-�#�R�PG�Ph!��?���������u�y���y��k��~fZ���<�3�kr���T��l;��o��ߏ��Ղ�������0�枚˙F�O_�U� x�V��RV�	.6/9�	>�G�IJZ�@��xɋ��o�u��3��sѬf�?a�����^!�����	׃���ij���U�x�C���9oE?y��*�0l�t��/7���Q`ᓮ{>��d}Xe^DI�a3$���dZ~�:FY�#�W�/���나P�[����4��#_r��N��S[���%-��[��%�o=�{��?m��9���ϐ$Y�G���{���;�������7�+N慞)�����)����c���p����D���GC+׮�{�ҵk0��6E+�b.b��Cs5/~$��[,d�C/v������k��}W�k����ۖ�R�:��s�������*z�}�^B�IFY(�F]?�n�rt����O.���0[�ߦJ���mlh�˺<==<W���(�꡸@�U�菋7_b~"��6�RG������$\��+��~Z�IT���I�T|����<>O$w23�s�, H0l�Ѩn�A�Ӥ�sqr�}41�:X�+6��G̷��޵.�"u���6M�z�bbu�E�n���ih,���>!���ϗ\v�065�-������}�����5;"�Xk�jr�__LMҜ.R�r�|�s#�H�<s����n[�+8�� �yp%�p��Ƒ+�J��K�#�:r��������lB�˺�;s?8����	��<��҃׭(��~,ή05���D�.�s�� 8�X�_��Xtf+>���ߴ��G�
����_��;�z��Y��	�(�G��T���F-����)��]�&:r�����p��j����@�����2w�-#��ѭ���.���5###f�����k>�_!W��K-U;��3`�~��#�_��|Ω�':8,C�

6@���E��R>�[��f�9V��Q?��adj��7L�[[gc�r��f�_�2���O��5����P�����毚���/�6��u���=���Ϫ���FjEDD�����0���NP[��� ���r�y�,�����.����b4\�|�l�3���;fo������4��l�k�wo�<GG�)��l$<���?��9�
y��@IR�������߇r'�����gՍ�����\Z�J�Pk���0��nnYR	��$6AN���~�Q�
����u;���]01Ȕ�n��D�7�WR��&=R���m����|�Eꍐ��DB
�0A1���w%�
�*{���H'B<�=<��㋄��Y� �w�}�$����;�\
Cd�Y�[X�||.4�I��d;��m�����r��Z�	)�!�eʆ �x�G��Ā�Ʋ�FT?� I��ם���1�շdZd�<8���م��ѐ���	�˚;�y�����7A��f'������/p����>����ꁘ�����J���LW8/��EQ� ���o߾v���D��4Z(���V�`�R"I�~��_�1�����Ɯ}率K��v��+�ظq��o�}؆UH�M�ɑ�\���Sʁ���:�N��C��g�8�[b�ns�˚4�`�˗{ �H�ϒ� 'w�8�|sG�]>>�$%�֯$�g���i@�?�c���Q�Q�D�qX\�����m���@3�ED�	'l�ܖiII���� 'e#G��ڙ�����GMì�~�{]�,���+���L������\}�w;�����x8N�%�dU��]���Z��3<�			Y҉A��,c���J�>;�{�)|��A«�p��R���o�[�'n�raQ�8'��K����J���V�wy�'�َ�_�*4ݻ��fZ[W�w��(�~�r�����j�A8 �8��V�	~l/<�ui���f�����/����˖�kη��x���gq��#���TY<��b�������\ s`Z����Q��`do��9�/�A�Wo]i��S��*t���*�.����gϟ�|mN �8�����1��������c��LDm���U�.:�D+�����uu��6O�)a�#����a�X��� Rx"T�
y��	ϴ�XS���6���Rk�s�yc9hm=:*i�
!�@xq�������|;����g|�㟜����#7�����Aj!��D��l���9���{���4��:��,8�1�	���zg�;Qc�?67nm�ȫ,��_��U��c�`z�azix�+/�	�t��! Bۥ��J�*�~�T0n��u�~-�ɐ����J�b�iچ@�m�sihmy�|6o���u���E���ʩ%��+�n�1[J|�
�u��*\v���_fuD�8�^��K�46�cW��:�2w�#�����;@k���"��>���;w�Z��ܧ%�B2>��7��M�W�޹��wA�elf�}���\�!�u���#vg7� >ڛ�L˵�$'!ʹU�b�*�N��� ��e�#o]�����+�:�<��'�<��8�v�|�~�j
z�%��� }��/���]����U�Dc}���oQ3���>������.��z���U]g��Y|��E[�e*H��>�Ƈ�ԑ�]�l�Q�>8	:s�|�O��I����~�q�����n򠾎�a�+XT~��'kAjj�*S�л�[��7�u.��J�һ0Ѯ0���<2�⣼�$ �h�����4�Ʋ��<R���1`㕕�w��%OX���������?K������ �/���k��z}ĭ�l��qV���;�*�Sς�j��t"Z�ќӾ�m��� �������#���J.8�������\��odt9��c˖-w��[�����!77ܠ�c&�UC^Y���葿��^齺�DR �~��-����6���L�V�A}�ͭ��*�>|�xhr�ם�,rwVx8�IQGWy������]�bϧ��q*F����QL������CA�v*Y�9�;w�v~~�jy;XS�������	��1V!�;�F����V��^\*��@Bn,��o�"�uiH��\V6��ikk�U����1ɹ�=�P�U���ǻƳ�4f,�	(���3[ݓ:�s��i��	| Jc��ywn߮V�[�:��K��O��|�X�h�Ft?Y���Ĥ4N���y�֌�#�0�S��?
0quu}~��V���Դ�H�W��W�%j"���I���o���|>�tr$;���f;�4���B�DUU�+[�$nܿ�8�H�:��pb<��H	�qrUD2�����O/�[�f)mؐ���*A�;7on��/�����9��L�������M뙳�{+d}����ǊO���+��L�򙚘�R� d������/G��a�7����(������6_Ȇ%��ԜZ2>%��r��A�����2Ѫ<^����l��n<�<���������{V�6�|���Z��Q�%������j���e%m?�;'g�}]�}�ߚ��ys)(%=7��!8���s�'h�N������l�`6�:�q/�էDd?��?Tv���ݻ�G� �W���fw�3�t2�����d}���Kw��	�?̴���?�����k���oK|�!�^�v--.Nt@�VQ�e�Ye�%"����L.,4el��d�fC.���Чh�����L�nMN��Ȫy���߿L�ulP�o�����K����3��O^M��O}�o�2��K����̋�	�&D���kK�o�4���eN��
[p-���M���A�� `���ANsi�r�<l��4ѽ��*�{����k�e�'����ۮ��ד�w�����|}Uל\\�$�qpH��'����/�w�����hbgle������'q� j�AII�w/j�� ���e`�u���6����SQQq'=R�b����7SQ�����	�5��f��~�u�4p]�9)��ش헥��ʖ��~����YS��6�7�����ϱ��2��w�j���in�HJ������`H�����$<��(���|w�K�'��_`���kͥ�0C/�x����C-�d���b���q`sCÍK��ܼ��ug����������g�i �1�!���H�Qx<���9�!c�;������`]"%׳��/^��d�	����[=����/5��B�����o����;�����2g�rI����><�����g�r�����e�VJ-�o����@��Q��c7|8(U�E�>��K��8�X[gǫ������塀�����f��m�%�ȃ��Pu5*��o�}�L`,��o=LJZ��ڊF�|�����I�5�#�!We�RZ?�>M�tUwk��Ϡ-eH�1����+R� ȃ7�⮂z��h�"A_�pA{��pE�ɹP5Øne��[r�j�����'�օ��)g�E��p���[���K6�[�]Zj0h+��u�2D���K��\��耬R�?��N.A�\ED����bbc�8�L��Ib�ǿbժZU�54�?���=�,��$�q�W��	r@�m�)ɋQQ�ǎ1ÓkTY�;�&�����}��SU֢e����0��<�4�z�W��ADt��O�̿.���,����/g>u�.�q��dWГa��OODh+�=1�"�_2���ᑃW�q�瀢� ��[���`�#4b�!i��xzz�v==�ւE�?� ϓ4�9wm���f\�;%�&O1��E�D�܌��GYoW�9 +Y��Ջ� D�Ǝ��*�����ھ8u�FU�B��̭���Ϟ=362JvnJ5s,��$���de�G��R� /Z���m�D^m����-s�	<]�k$����5ı����i��F.M߰u�E�3fy驩�)))xBə�d��9h�!��������̢��b�u,�d*b����f�҅����Up��tnTlr� ,�ML�b���ۼT��#�<n
�x~]�e�N�5k���Ӌ ��7R��b��V�~�������"b�5�IL_g'']���vo�~u��z2�H$������TTT<�L����m�S2������7y��<6+D�]��@�3ٶ�$�q7O�)��<��u��q�j�+�s�?ʆ�Ĩ����w"����EڒP�P��ލ��X|o���9E��L�H��@��,�K|���K�w��?m!߱..B�R �Eݭׯ_��z�~�
�r��I�xR������p�ӈ<E_����08�k<u��K���F��r���t9IP�=Eu���7X 
�Cʻ�?�̑�������y�Gw�cy�g������[UK'N����Ͷ	�(`Ïϟ��i1-���ҷ(t313�ο��6�Fs�q�v�2�8L�V9�+Ʌ����_�ƁO=y�y��{ZW�^%ώ���9�	a�᲻{1y zVƖ�;�h���׫W�RS��V�r8��ڮ~����������ny�֙IK�X>��6����?";v�(�4� ��d)%ʭ�8X!��̥�B��?oߚc%K0-,�R�d�
��ۜh�]^�5`��x6��$��]w��E���RJ᧊t}�y��R���u)�ғφ���������D��b�Tb}h�C���`�-���xYڠ@��Mg�ˑTކw�&�3���vH���k�e �E��;|�i@��׀)"��$��ϫ���\�� �m��'d�xpZ!rsVi����]�G�W�̲e�/�Ф�����׭���a��q�	d�O�C2K�B�°BC�<w�&a34Vœ��"&�0�Z���\,� �=�g_��f>�,�p�Y�PɮY��n�FFgH*���X�\��o���E���G�JnV6���d��ITrK~6GFFa�}�r�����!���\Z9����,,,o�d���FC`VW�\!O�u�Z"�?�\<�$%�;������H;��l"������?u�aA��b�/^p�G�A�� M7�ڌƂ40�/�W�Us
�W���<�=u{���OXy&�3eٵ5���͂(���4Enɴi�2�	��Z�����==N�t���g��Z�ǅi�I���rk F
���;�
%�>-�]Y����`�J~a�E/AY��Qܘ'g��Bۜ��X�����5�,<-Ԥ��A�T����HE�����5Y딕oi+̀���� ��I5]���+B�iw��'�1�=�.Ϻ&���hXg���g�n���y,��7�I������2�U BCZ�����nU�#�R�mʘ�MA�kq��Q>�[�K��a�S!.��򗭯mij*�b��sf�ׯoWVj��� �|������F��qk�	PGk�EN�����\�
�@s HO��L���hl������M�]k��������P,�(e�2>��C�28]�@���b��2��7�<0���rN�<���Y���>>>�(��
�!G��C<�Seպ408���g���e$��gWF�~[��P��y��ё�+��Ő��{���(=9�B�/}�a�����Ԕ!���D؀�z�,�nޢ�����o�ۏ[y���@��٦t6�����
���Bƍ8�бS�[2\_��[_�!: I��c˳n��'Z�� �1��QrO ��6,��o[��,��]��ѣ6"�����W@`�4Uǣᐴ7��W���pOv?>��Ԋ���KT�,F��E1�j(x�U<Z�Қ�|�K��v]L�z���O1�*o�8}����]o�n�0V"�'��B��W$�x� ���
[DeC��k`K+�s6F���~h�;���0bH��CLv�l�ڟA~�@n���C���zc�N�B���ooAp����ת�� �C��J\�0;���W�1�n=�=��b/<� ,fd�|���}-f�h�,���QB*oE�������lr�^p��9��ɉ��!!�DY�Ǐtď�b�t+��j�X�=� < o��X\y3�������*Տ̧�s�6 	*d��m���ԃÎ�ơ��^��Z��E���ڀ�{���OD�V>��}�ˀW>�����9ŏ���;��-����?0�pݬ=�������ON���̿}�Ύ�ܝZXh21`]|�Ӧ��w��'�����zEE�c,Ny�`�ʌ�D�km>����͛7�F�������<�ܲ A�m���[�GL��:�!'\Pa��x��$9rY��Ǐ�̥�R�]�����H���x~8�8�����	&�&��ǿ�9m�nĕk�/+�q*^W���X���?�f�Q���#,$�G[����.����ߗ���x��� �l�:M�<���6$M=!"*�
|�?G2,�.L��	~�W\��#��Sz�L~]#Q12:z1&D�f�+c����m����ݖ��P�N����e��A�x��9r�ѣGQ����7�����!��� ��'!w����|�E�����),�OXke�eKy��z&�ޯ����)a����9��^c���>^j�03�~�����Y�Z�u�l�w.ã�<�ٌؙ>��X�lYuA\�'�r�.#��$�5���������̡Y\�����ލ�g ���� /�2utrbN���2��,�
��y��
�qtt�Cv�����'zS����p�O�h=]a�!��o]'����:_C�4�P�R�v@&݀VM���۠ڐ]ɛ���ޝC���e,�N��N.9��1>����x�(��9Q.�k�B?�m窔�#�dN�W����Ct̗޺m�ggƸ�I҃�W��cR]����Y����|�6�c*��M.8._W������%KT�75>	
�?�iR��l�uy��j_㇂��
Gww���V��_�Sg�'��&����0Ǆ���fkx��y�t�O�V���{��c��_�{�Gz'>�hzz��l��,m4}�@�S:�Is���~�]q�?/�A�E�)���J��}�O�##��Iˈ��ѹ�lm�b�~�C��{_��J|���9c+Z��%�i��2�{ڃ������X����`B��TI�DV�5�u��IB�E�����x�~~�J(2���6Ѥ9a�]ݱ47]��)\��Pk #` [�[��m��X�sj�g7���&����/�����/�Z+Y|���<e������S�X�Z���H�W�<��D,}�?]��BԘM���!�ZQ���|+�b���j?�d������H�Bk9-?'�9�������A�)�i;�V9�4�g��QOu��Dk`���?�S���a��^�|)(.~; EٛNkN�`�_���A�Xק��Goc�CL����u���sm�������Z\�e�ݿ����`���X�ï;;�s�lx
N�yf���_e���Oה֯���-�
d�������� �0L"2����ã�Ѷ�X�뻡`%l�����p���*,���ӏS>@�ߢ@� eQw���i%��,�2�a���Ԛ�~���q�w�K�v``�8�A�W��SwRۑ���<��to�av}J؛��2���S�/�!�v#􌤙,�o����1�TG�J���[s��4r$�N���_�C�b�)fMg���^)P��H�'��3gμ�Kh�8ƨ2B�a"�\��q�RҤEq9 N��Thm��e!�|����Z��^S/�lw�f�9ƃ"*�`��ttt�p�\bx!۠�*��g���?c�|MP/|��G$���g#ӵ
�w�Oj�k��⍱����L��ze<���\Ƭ�E�k�A�arH���;�0�i����Jh�qQU3�=˨\8�i�$}���Y&��^"����$o�����=�j%�qH1�`o5��|�k��^�>uU�̯*e��R��1�VvEU뤞cL"e�{%�&�~�)�C8>{�g`&l ���5I�i�Dԙ��?2�'{d�w�~�p��b�rFk�l�	Z��xç������a<U(n*�o$M�+>��1�Y��E��
�������+��d2��`sxC�Ŗ�xC䎔K�Ҹ����5�.�C�N�! ̍Т�B�c�A�l$,�,��$�kAK,�Ԉ:_h�y�I	�ʒ]s�@�rӜ����+�LYմ�v�D�W7�� -U^���K���"8���tV��"N���rD����_�`w0݄�V:�o������2��;	j�`+�ǵ�+8����c�/YZ���rB��Z�K�~���lD\kK?6jR��k����+=f-�6���JX
4p�?~�������6t}7�\&��� ��y��t���U�u�����? ���*���c�W��v�^R����*��=���c�ب{��;����b.ChNl-��ݔ�j��f�y&�YTJ<�
v��݁�{��3*� ��'s/���$_Vq����O�J(��X�OIS�8�����L�̌ցt��fc�IA�"m:^6�(�ƎrbA,̚�č�uww���`�噱;v<����bߵ�)uԌu�ηč��;�_he8�"δ|f�ɋ�f����R����O,��b��F�ϬQ���O�$ު�`����w+�SZi�&("�t�g����GP6j���q�ꆏ����U�!0J��Э�:� F2�Ak@XPPwz˷��al1�3�d����{U����*�|�yl�ڋ'�}��,��̽�V�iӇ���<����P�+!� *>!!aŵZ��죔C֫��"�g���se}�,y`2ҵ�����♈繬��ò߉|�z�I[�*e0��!�ρl�����#�x��9���Ǝ��Z���%�i0i| ڕ���gdx9I��Z	E~��Z43�n%k��M��+ ^��9i�)��0���/��7Nb��0gAmijk�~�05xh�J����ʊ u�O �H�1�	=`�~��4W�:� ��Ev%{�7��f�q]k*�m@` �<�:ᒃ<d�Y�$Bn������y��'�����-^�v��j����iXrk��e��=��
�k_kA�� �mDg���Ֆ���T���Q���szPU�P̫nn7�����j�� $:se�LO,|۫�p�4Y9J���e�5�ˮ�=�t��qF�LWc=Ǿ�Rt��k�[::��	�!���	�2�s�f���zHVn�Q ؙ�r��(�<�c��=���,��		��A�,Y��bG��=?<��b=g�;�"��I+��vދg&2Ņ��LZ�>��:h���R�T�5��ʎ����9�Zq�:{oFL���Q��kK����G|[U��3����'�V�E��^o��]�yA����%��ep���~���5�"w&�xn��BEM�*++��*���++�t���>���V
[�����hG}N� �Vj�����s��s��/�z��j�ÇeQ~z3�MßBBBH�Q�aXB�(D�|���O��fDb����[?O��f�w�t)0�mϋ�V�ӊ�kxѓ���H�jg���2_H�!,"��c�e�Z[ooE�v^_�g�Y�T3�2}�:|7v��3��@^�����=�v��L~Fp�nan;��CCC�߸���p�m�ņ�Xu�׊	5y�dZ\�Q�ˀz�>4r'Y� w�0���3)���G�	�/�w���[����@��C�5,��Y����&@��z *˴�/~��y׌�v�2�:�`%4=
!�n����*B1�g�e�/Tg��B������Z�`/mpk����[�2��G�P��B �~�h~x���S$W���p��niQrĕ�����x��`;v�	�����C�3 �;���.�"���'ѠNV1�&l˱����{��9�^gpd��n�
x�	v�gcg���};��w��ࣤr�\��<U [��qq��a,�����a5u�ŦB���8����f�6�L��s���
��7��2��71�N;ԝ�?bk�Hql���X����ʈ�6��z��1'D���;�V[ j�A���ͳ�|{��`t,����l��c��y�dD!�Hp�������f�n�� �/ 
����b�NZ�n3�l�Ś���euQ�e�h��(a�� E�Xy��5̀}���P���B��c{�����'�	`�T�8$�?�c#�S\a`��5vAA�@��Ǿm��a&��1�م�J0C��K�9ۻX�c��H�ӟF���&B1
���n�ʳ��c���J'��B����GRٺhZ��:~��)�
�]�v�3R�ՙ`u�m3V�x����H9,�k��5Z�FZ,�a5���dBA6g�.��
�#Y�[�}^�q��:���r��)'!��������������h,܊�Ϝp����#Ǿ6
����� �+��mutt�F��8���
��3N�f��Ԩe�>���J6Lr�s_���M�'�Q�2W�73��P.NNl�����V���?'��m�"T^^����P�XvycE�ɪ����Su�Ũt�D�`�&^��+�Z�m�\FPo�&qU��xFб�_=ܟ6�`T����us�l��6Fm����𺀾xx÷]ha��?ݓ�̫�n���׶��`����Y�8�aI����ྰ���4[q��W���mٙ!O	[��N�FZ�v�e81�����Y��1ܻ�^��r�����S��p)l�3+���dyE�+p����w%���U��e

��p��S��l�f>l��	+�Y��R�"��:!�F�)�k���:)Ǳ���������m�j�m�J��l&"�>M��}�7


�9$H�:�P�0Ya�S�	mq�E�v&� ���h­�z�X�j�n$�H�	 v2V�D"Jjj{��5�gī���Q[��K��	�w�bo�>Lb�����`���-+�$��ͪ��zS�-�?��FivNN+๊�؁�FӚ[�v�;+ 0<8�B��=aIm��_�JN;����:��h��Q�'#D��ɐ��&&O��hT����tEEE^P$JX 9\dL;M�Kd���K���1pF+r[�#���-w�x��M<S@��j���Ә!}U@7�:8)��4�b7�(����h-� >�	����qk�oΰ;xP҇Mq`d�K�]�^y��x�����HL8�Cv]	Ђ�i�s+�A�A��@�1�n�2�<�(�ܵ�e)j�ۇZ#G�r�D�r��-"���s��It��֩�
3X�g�uWyn$	��-t�f���>�$�\8c��~�������]Re>��~+))	{�!��߀Φ#*cl��=}���6WVc�� ��zʎ��DO
;�Y�oӶ����^�0�3����\�|�5�_	5P8������#�z.��g�C*~��Q�?�O���z�G6>�j�bK����B;ʽ��j@��A���:���wz�Z�0x�౮CT�vtt�ąr�؛\�) o�'l��
���[ɗ�}��ϨU�iǣ@�{	`�
Vl�	��AV-�qr3vnę3yY��O�3�-H����w�X vU=��j�	Uە�6	��D�$N�H�՗��9�a�i\� H. �,  �)��F3�s���&̟a��֬��7ia׆-��w� ���ᪧ-v�255��&���1:�G�V�����ؘn0�������(�t�]`H���y�&Ҭ�E_�~�Ƃ��틲��oJ� �[R�b�GY�����ts�����oǦ�e"s�>+�9Q�f����23�!�J;BJL	�i��s�:��O�GV3��2��`$�r���*�p+�T�еȥB�KԚ��d����x�!�`j������!�1�
�>0,/�1��896ޫ)~�X�ts��������lق��Ţ�$S�2��=fv�����h�M� ��p��1�M=�4Y	�WX����㕭h����#��:2:px�k����o< �E�&ȭ��dLz50��72*D�W�+�H'z7�O��E!�׮i),�b���|ћ��%Nd�(�X�N;	~�_����뜕����1p���se������ p��h�އ�v����|�+\zޖ�oW<�^-��D���M�H[?��f�j0�zS�~��j�� rlu)��%,B��='����ַA���3�B�Ug����?��9����g����I4'�+	�ɣG�<����y����K�������1֘xm�w��_p��ޓ�w��h� � M�¾�I k��l�VN��� ;����	���y�=���f��MMN�+H(�ps��ϟ�c��u���h�1�1$�"���Ò�3S�C��<�b���������ua�	�cJ���t���ߐ��ERHHֻ����̹}�������3G�?oq�qf��@�1H����q}�z·�)�f�8�^i/��`:6��U���-5�6��&�/���X8ۓ6���X�ct�f1�-ja��%%�w�=ִH*����uv6B4���L:d`F=}cA��	~���$����u;��,Ì��pw◥����5�m�g���`R��NΜ�����dQ��(al�c�]��y��ͫ��g8
���� mX3~=}�t��A/y9�HU���»Ӎ�b�Ep' rs-,�����Ƈ�Z[����%��vN��~����R�2������T⹨�	�����ۃ����z�!G٨��:|��,���0e�?�5E��΀�0��\�����y��11���1�g6bbD��-����d���0B�9h�o=�D�fv�Z���X�{��(��\kjs�����䛃PY��.����w�4���=���Z������([:�}<6��>������[�Ӵ��E���b�J��oP��$��Bü�R&�+^�޽{�>}��~��݃f���۞Ţ��1_��El�η3�%�}��+��"���tɕB"�{��tV�<g�s�;� �N��7��k�}�.읁�M1�ZI�<�������V�'��1�71�#� ay�Ϫ�132��`s���^/[Z JP� �D��s��@L��K��},�o���g39���j'���q!!�3�A`pաء��u�ò�,I�!�T^\���I�Ý!���o�r��X}�֍3Ww���(�D7s"��F�����[���#���ۀ��8�h�J�G��UL�HtF:�4"D�	�� ,�e�����\YlɊ��go�6���q�ĈpZ�s0TAHÆέr�56�	Wc�p�3�Ȼ<
�kc��ao)�O>l��,��g��e[��A�l����ӊg�}	�]P�<�Ӳ� �:��e���$�6�sr����IWά�9V��<0����z���åd�}`��އ'�f⪦-�����F��J�Uf-f;;�AV��|�u�aXƙ{�S�Y����z��f��"�X�Ǽ�`V�� ��:��^��b�!���b�i6�����cSv�#B�p�<8�mH��i�賰��5׌�-Lk�J���^����Q�9����ʊ�l�Ӂv�}�V�y���$'� �ʏ��(.l�bx&Y�����Ǻ°�i�5G ���ʿ��B����`_Zƽ��2��_�V��T��hF��ꂚG��t��ޕĮd`�ب�\:�>�xrrrү/��M�t��M��z�?o�!�f]U�Ob���0��߅A�������bj�w_�r���Ǚ�̫�@� �֊��K�ut�O
X�&�m�' q�&E��ܩ��P���^s�!+{�p�ģ8X�̜���6�3����2���@'d�>�#�9՚J���{�d[�]����gk8'�1@H�!<�Z,�#�Q �i�q�/z�����ζ�h��|�x��V)\w�a�2�y�=���X��b��ꆆ�$4ҍaTJ `s�?��<�
�{1�����G����x��C��{���y̆���/px��Uk����ث��z�77fgY9Դ{��E+�[a_��(��khL>��fu�V���_�o�0�������C?��G��4J���(M�⺂�Ʒ�Ko�{��gZ����"�:ܲ�Y]�Rg/��bUY��\�Y�?�T�_�����iuLN�Ǐ� W�ip��y�)i��gx������`؛<��}M�**BxԨ��F��o�85�5�N[[��O4��*�2�C���L%�ōWg����11>��ގG����/��~��^4&�RP�9~5"�Z��&��e�Eك'�^��m� �>P��_���9rD�>�м��7/djOˁʹ�NK��W��*}�n}
V߽��׎��S㣅�z�,��h�8fH��>bӠ?�S�O�&`��zj������\o����nę3g�G��׷�RjU���l?��.-��qr/���(� G
S�_X���\�Htl
X�Ǻ����"�=w����0�;{J�n
j���x�\���
�2@Ew��ġ�/.��X�.݋0�kL����e��7o�#��<؛[��M���N��?�ǫ��yvt\���3��|�"�8��L�|��t�@xż�)�޺'s�]]��<�
;����� �h�%��rMUa��+��+���=٭ ɦ��c�;::�F�M�]���?i���V>����B���t��	���vUҏS^X�������� z����Z��[����x<�Ss�t¿� ��>p�Õ�����q?d��S���u�+�؁��+l�'���j�s�ʖ���=��I7�
��z����{R��"���>�!2Pd���HYq�⏄c�N��Q�kş�RqD<��ӧ'�Tk�4���.EW�sZ���-�>�a�� �p@"�<�# ސ���޺���,Z[qG�*�/��O�/`��?x��5��i�c/Nn-�w�0b���~��@��!���q����3 �x�u׮]A=[]�.t$�=�3hb	fb���<,��v���|@1:*��+[�x�>�l�6�
��w���^��Gz�m}
�*��@�)�t;j��w���G�Ѩ�@w��$�$��ȥ#�������@E"~v�h��=�z|�+ׯQ�Sʒ����!��ޛ����Ii�b�yĞ���,���X�k����!W������N�gO��ѽ4B�6f��d�$SO�+T*���;֩=E��[vD���Z���L�Q"�!_�x�/�Y�w���Ɨ�w�i�Q���W�~�J��C19���Q^��ٱ&͉&e���@��o�!��ʔ��e��
"�YH;��H����@K�6�\�|Y~������	։��⢢�z��ކ=�������̟,�m_�]�7'E�;�R�>�*�/�Rw(k�x��߿�G�UVV�����
o�7-=[�0����py���c��F�>H��X���hZ���ʿC��'��MX_P�R����z25�g���J��"7,9@��G��AQ[[�����x�l�hS��]��J��o�@��!P�79Ih8u�'*8�CN�ih���)����p��C��4�v&Sl���=��8nȼZ���R��7&ዀ�!��=>�)�L��J�R�y~�O�T�o��t�џ�H�xI��y9���x/�`�V��3�!M���gv<��N��U�����
��m�U!�:����j�>W��9gqK��ʹ>��˅����q������\�m�ǰ������v�������C��)��+1�$�cw/�;9k��� ��~�냶�Gھ��{3P����)�oT7�U������Z���6h<�i��%���d��ǚ~�G8���+p
^�.��3�ߪ�b�������7�zh�=\�c��={�<P=Y~��Y��q�6��2R)���D��8��Zc��>^��#bu��}���fY�C^�����{q0BK���'�C���$��}xp]zW�.NN'oo�}�ҍw���P�����mjo�������6�����/�Ic3��;wd2��3=��L.���CP�W��;&�|��X�$Q�����w�Ը��k�b�v�̡�CN�3�Ni&��
�,D%އ�L��w%)�
e���S�^<�BQM-��I���ķ�뮿z�:ܽ|���e�d��Vel��FAN�5x3GS��@�����;$�zA:}���O֓��8�*�?E�ˍ�u����7�����!������� �޾�q�\#��d�����o�I�{^�x��rM���P/e�T�,jyb}Zc�!$��9���I�l��0ܼ{�[�������h9�ʁ��G!M��V�K#��ŉ�H:'G Y����6P�zB,�|%.Ж�\�?4�J�� Y���|p���1cu���ʢ�ᇅkך=��`@��g�AOOC�_5�rr6 ��({��m���)4o�l9m1�V,I8:j����E].��6�� ���C �A 8��P����e��W^�QS���L[|�~��=E��H	��φ1u�o�2W��C���x��x���X���D�� ��� `� �@�z�Kk��d�.2QQq
�Trko�w����_���(�V�D���~�F`��͇2�T�G�ȶ���}��.��̒��6M��O��=�Ѵ���e�%v�\���4����*��M�\6x��C���ܬ.�!��{f���oޘ%������XZ�G��L�G�b��q)<�+�NMM�US�k�{�Ň� T�-�<�GZMfϺ�p�OYA�~vͱ��o��Pm~}���{�+�z*,�/����{�/��9����\sBΝ���dne���Շ m��{-7wh���,*���܍����s���ۼ�4��Ws���o{|d����c�N=R�f˅#�\��jdd4���oP��[E����o�(�K�Y>�<��ĥWw�a�2��|��d=�իW�=���M �k߆��Vbk�E����/�o`9w'E���ΫL��[S!��n�0c�F�
M��@Ugx��v�k�?C�#�t4/��\�
$-�1��l�R��6�o��b)ؽ�V�#���ۚm������
b>�}��<
7��TZ��ԇ%r||�cbb���<y\-611��M}pjN�<���(w�s�$�P?�ɛ�*
�E��Z:�a�O_�r�l�:v<JK�1�`��
lnmM{�rϋ�ϫ���e�c�z�݋NQ��o�1�؛���e��w�#�;8:�hN}�<���9�8ٗ���<��o
2�	�|�W���D��Հ6���@ �c�����哓�.������D��gVev�(��{�\|V[���RS��-��e�үk;ӛb���&�/7g�`?0�� ��'��6aϽ��։�������Z˗/OŕS�򋻤|F�MFFF�mm7���3��3���Ibu�
�ۯ ��.f��͹��#Oߺ�����,]I[��`��5��n� ������].>y�~��T枟F⇂tJ|�6��P��.��+�k����k�^9r���{i]���~�"���\Ǔ���1�>����p��E[�43���Hi|�*����A�azS�LV�%W#�+ tJJ��_zS�'D�܊�E���r��bq�;w��ǽ߾}����R?P>>�1���a�.m���x"+3h�~�n!����ڵ���^�&��� ;��/�~�d�~x�(l"u�l���#���|�R�klhx|K����C?E��B�w��7e�����ޠc��M�4j:�i� ��� ��$5?   !���нշ��~�㛚0���P��~|>"��WH ����=����u�m_�`d������X�v�<W��-�~��/�&Bb;��Fl�g�w/�;�P����~�
���δ�����ڌ�/ޙ��?8���=�M޷�/)2KypS?��s�m	.��������U��oѪ-[��V���pD�}i�1PO½�U�S,���s��X�m�֏�@/�c���K1����F��y���Jv�x�[�-Փ��ӬT�7�����v��I�}l3��G#QV���}8Nh[�9D<���((h�(�L�-֪���oT�WO���_}�o�H� wT$Q���~~�j���"~u�qm�t�~�:�F�������;��6<�����lx�U��tYi_�@l��=�reAs j*��.ޟh^�{'��'��7���q��)[�bU	��(wۗ�5�4�nQ�8qJG��W�үg��A%&��+�������C�N|�+0�Q�_Ɓ�E���������mZ*����+=9[p�U��s�<��,8	k4�۷o�cr����zn������~�"0�݆=<��9Xm�c�TC�̓T;��ي`gh�l�v��IIe�o�ؾC�2�/kI�3sW��F�/RI꼴>���!���ǏV�0�&?z��p ����f7����b�
[��j&6������
�[5��1����?�5���QҔٵ��X�ʓl�l���{��K;����%0ln��r]�0lA�_�����g��aٌ�V�֋�t�������V��~�b���/Gb�0i1�xt�RUS[��~���ڬ�l��.Q�d ����2'�kP9+l6n܈�3דU��R�˿��u_�+&"ף�-�-[���5,@�N��(�޹>a�o��5;�൴�lc�L @�S�[N�:��8�EP�!,]�Y�*�@9�X}fh��~d^v�贝*�V�2DWY	fXX�_b�u �wC����]'�2�:qH�AL�(�3�ZP�xb�I�9��<�'�*��̅!�����dSC���]� t�=&&)CA�j�\]I�~6T�z�
X��(l? �x�9��8H�*y}W����}}{d��^M
	*"mx/$V������N5s��(���C?4y�oL�hvr��ց���Y:b�[�\��0$d��k���`�.�8w.���"�]���6�f#� ��򐈄���IH��g���+h[��r;%e�cmZ��%	!��X�@���9P���.����M�m��ނ����~4*<�-U��P�ņT�X�7��t�K���R�<��kc܌;����c�;��L�nX�U�	J4�dQ� eH��"9)93�"�JIr���$�Y@�9���'����ǳ�Qf����n�[]]Mـ��p�坽�0H�jۧ�=&��휁�#@
��Dn��Y[ZBq{�a�fg�w��δ&���}���a���H_��j xm���JJ��[+P���������/
�j��fh�b�U��+�*U��?v��6����+Xmym��?){�ȵ �4���F���9����U�!]R�m'T�Wl	_
&�+U��y���N|���=�9��>���f1�kN��`�����I��W/�g"�xh#c�w�H!��]��Nyyy��i{g�'x�i1 ���]oϡ^\?_%����U�N��`��j4��U���/'�:�������`Eݰ�ź!��w��gK~��y�
���b��U�����ͥh`��]��G�_�Y@��	�`�.e 5�����x�)�B�Af|�0T@�F�nA6����r�%��� :8}4a�0b �e 6|����2�I�9N��J��E_\�������|Ϯ$/J�z?�J�� ?�J�ؔ+ @ި
<�lL����뱿(a#m���[{��{���˲���v|Y�� V����Q���}o�e������ 0C�����ǏM
��d�z����g�GPكs��)����\���E�������|	�s�y{Պ]�[���Z{z�C�v>@D��eHp_mmmD�C�����w��6�MOW|/n�ng�#���y���t~��:���2������N�@R��Pel���k��iUxG�S<�q�R�2�nDd���>yBaT��:���}y��ki;�J��cכ믣��p$�S����F��Ҟ��iMM�Ʉ �9t�]iQ���:�/����uE"���*�F��0��9#��ϟ?aC@���8��g-U�'���g��:���n�I/b@� �3�:vI�[���|�UFc!lO&�����4B ��BqدJ'=���p<�1�齄�P��~�/R���{��6*q��!���
i&��%��LNN���%�7������k�G�P0�a�|��q��)P�9|������@W3���)A%j3�S�JP6��i�N��.��8�~��;^:�y^h��~��HB�C.X1�C�i�����2��� ��ځZXc�[bN�� ���).�������Tٽ� �F�JެP>���iH�����6g(������vnT�@6C��<*ג�3�E"��4�&��I�8��N���-J �rO[;rh��Zg����g�4���^}|#�q!�8\��^LB�����#�������˗�QB�'���z��Z++,�A��&�QS�_vP!+G�vg�7� B����Y�j���=z�Cv"M�VW�?"3���}6�<�/^�B	

B�70�)������(���1�����֚o���a!hX���@Y�77�T\z���M���P�1�40�	��KJbQQBX�� ������HZ���F.VQ=���.&	
</�êCR���`�=�&�}}|!�� ����|ow�9�n>��C�*4W ,���dj��&����� !�h߉������G�,L�z�v}�B�c������[)�䴰�_��a �C,,,J��-āW�+�S&�����g�߸���5�u��cx���;������
�K��q���
,�e�r�<(����.� �x=!/������~�CgExo�t�Tո. �a�0�	@�fg}�-�30R9S @�����d��)��Wƕ;�֝$um��i���W�~�������~���>�}�"d��e!�s´���yN�����e��C���$����d	`>��ɨ�Dc���}||�߁���)*I";�0�����L�"��zDRw�.G���@5@Zα������QUh���C��/�F����oW�TÎa��Xd$!�y%�H��7��6��\����G�3�s'`{Z�K	f��N�� ��}� �z��������\u_���@���<H�ˮ��㳧�����.��uN]���� D�L]خ�اpf{m���˰�"���a2hJ�ӯU숣�DY���*���,~��^XЁ`�mt���@гk����*(�OP�����yRԢ����A��'�؈���� 
��z��8���M� /��"��PƐ�l�wmmm
�hR����I)�Q:�6	DR���,m#�XwC�}Pﰋ��zK�T���sG4����5 +o:X��a{��u OJ�����G~�ػ�N�		u�·�'�В���	,G���|��
-��_ ��l�u�����P �@̀��@J�������\t2Q�@��KT\��I�b2�,�]e��wuYW��8I�!�I
��A1,,,%���7>�R��na�Y:�F�;X�E0�`T�t�
�oÛ(���;�Q��u++Y[[kf�ק�Q����y�+ѯ3Ka/bW�.gZ�S�Q�b���Y�����,L�'�n�;:����5�����_r���q����� (]J�7l���$Vo��>���y�����I1�޵vvj^؜t����Ot���#�� �!1����$$FH@X7����v��"���'`+� *-�G���F�p���Ā�-D�����6M1b�bG d���C<��M~"��b�:;;��v@�������O�āG755��O�
 t���г��wDxxZq��z-��x��ߪ}0���>,�t���Tom�Ѩ+q&M�$������9m g �O��i������;����`�C:����|
P���|"�,������ ��_�|�����ݎc=��;�מ��\ȫ��Qg)���r������+*C/���t7d[�f����>Ϥk�X��}� ���<����]:�΅Ċ
������ِ#�'��陙�1E��X��2�q\]u���=���a_��A4Z�L�F��sڀ�Nt�1���~���<z���Ψ��En�SC灷�X�~�n(
b)B༯7���:��&\:hY�br'��L��5�yp��7�8�d�m�YW`��ɴ�

bW�8�X�Zs���x������?�u*�ב�k��<��h�R3����[0٭�BAF��&lv���l��X��.�/����ܡ���˿�P�ttTo��;�@�Ng����qη��� ��� ]
<X޻��E	�_�B��+L�@��y�K��$����%�Z �28�3S]�_�*�m�;vjdh�))� .��׌<&�@���)�vD�=��_�5B�;B%�9���<�[������~yy��Q�0�.|�lO[]�\\K��\
�+��
P��a.ܵ�Z��{?�܆|�*|�
}d:溓T,�-�AA���<��OX��RIE��크`в��R���-�&��bو�l��"��V����C²xxdπ ̰l���%���f���o�����Jc�s��?c|X��������(��cA4�ar����J����M4�ml!i��mӐ§:�ٯu���H��f�='���cR���Z���.Ow��#��:�B;~�WS������f���z��nʒM2��4G7�����%n"E��yy�d�c�Q$��� �P��}��G���������y]\]��Ђ �:?�)*�8�r?a�X��<K��fWN������g����)�<�F��*ĻթBB"�pKO!��㙙��.���ʤ�e��l�i(خ�����A���ߨԹ��Լw�>i�g��C�=|�����@�{�uw�Q:'K<G��	�/� R^��F�Pc���<�y��Y+��p��3�;)��Ϥ ���3�a���H@D�	0u�:�%ȝ��,滉7ˡɍ���Ȱ���#�BK�Pp�Ѻ@� 8�<�<�Ȟ4�frE�L�{R��p�&�@ �^������n&���%�������yy��*�n�7w.8��\������6
�j����kddT�`�v��y���a@A�7�c�VVm�M�	���o��x���7�F���~� Sw��Y�%��ж7qm��y����o�r`r{�,\����%
�V����c��2�E6[O�[m�.����?p�YH��< X��pq���A:H��O��Z�es�TX?�r a��x���A-Aף�����l'�v�w.7x"""Rޛ�@����ʀ�p��n���M�_8�R���D[�4%���L?�@)�K�$bIm1�"=M�u{g^���J�&E(��L�&�l�c���*kȘ葟v���D��@��m��F�(�%xP�r?�㼿��x�/2�	#�^|��ׯ'�6��77�	Ύؼ�~�3�m�r������骓VO��)V֎��ʬ�����Ux�a�����߁�]�'�B6q��$[-()����S�������h��,�����^���<"��o�ʌ��vX�/%9��˱3@"���tD
�ɓ�F�n�TNB7t'��P��{ L��/%�Z��ߑ^�؂������] {#��^�{X��\�Fx΍��J��f;	c0��x ��?�w��ϟ�a2|��`����yҺ��84�9#C� �I��۷W���VQ��V;r�d0� �È��[c��޸��VUa�n3]���D��I������֖@/�\4�K؆�S(�6��*�x�RC^�����D1��Pɀ83b� sss�2/ ��HA�w"�L����$@
X�F�`%�K?Xa+�J�JX�C��q��DpssC�TVV�&NM�@{x�VPP|43�^2�E���\(߀j����x�a?P�0�7��W�8�q�}��Pn��Ʀp���lⱍ�? ?�`B�\o�	!�(LI���խs��%�}/;��Xܰ4���-������\�P��b�.�FTF&n�U�
�L/��^jr��6���<z(G�A<<�_�,z�%�.3J�I�P��N �:��Ba���m&҅�ZzzV$�%sP=%%��ɶ$���p�27��U��&��0Q��x��VW����B�J0�23�@TE�`{��zmw���#� ���HK�����^CJ�+&��@�wi�ۂ��iiJ�(��D^BX8�%��˙��@�7;�S��#]jZ65X Gz��w�%��2���cv�U��M���__�g��T���6�� L�?";P��` ,���G��*�i�Gڒ�����qqp?���aA�S�ɟ�
UI��XlV�Z
q��uH����g0˫o`@H/ANL��p��=�a��#(0R�ٰ�`��T@!y��L�r����|�e'�ԫof�%����,�92b<��8���1`_t��񪦦� ����^<��Z���g�����wO�k-tc�K6����LtW�q�~eK�H!x9�%w�����&Y��nOG��Ȉ��B�H��F�l�_H>�� /�+�P��Y�P2Y��E(�(:DA%��R ��Qd`߂1*� �A(��e�q��_R�!9��!}�~���0l�
�Ɇ��ۋX��.a߳I߽o ��ȭ��=��m��-S��W��[Q|(�N�Lr�����1�(K{��Z��u����4�AQ3yI�Q�j��w�H�"yS-0Z(P9ЅK�|[���A%�>����R�wkO~٣|y�l��g���Ծ���t�`Z/�cկ=��U���������W\a�<�qp��a�����Ty�ޱ��Ur����G�b^�2���ֹ��O���^	ȸR;�} �p�W�V򨯐G�
h9�wu���,�z�,p�#�+��lTu¹8��jj	&j~o��P02oi�^R�Z��չ7t)+�G���š��Ñf�:�QYu~���n�8�]3a.v�UGZ&���������k�@����*�x
}���@\��z^*_�����4*	QϠg�c�_R�X�L�85�϶,%�!P&���R8�'��u�ЫW�Ǚ�O�h�;s&?�3)�j��֫Wc����ǘ��n�_Y"٤�:�R���#�L�HY�����\T��cv`���
�:��<J�<���ϟ&���y�h����;@O�w�;���n*��JS�qF�P?ф��c5?��?J8:z�N�4b��u����N̨�JI5���G�X^e��˧񛚚�#a1�)�8VDv~h�'x���#r��<��H��NZH�pce�`�k��ꨓ�r� cɇ�L[������� 3d��y����������Ⱥ��6:!w�e?������\�+,�[��K/�~$j�pp�<�)��
@�2�cϨ�`"�Zb@��o�9jhl7�c��>�����e'� Q��������|����2ñd.@�h#�8����<~�D�Ƿ��V�5ӧ�����ob�=��{A�*��W��^�-��VTF��gs-�K@���ʩ����Hy�<�+ѝ ��e8�E6ڀ2�����N{h|zC�-��z��Pz� E-6���3b���gu�Nǰhuwz�٠)	Ơ��dm��������:j����Ð�I���U�|!�H�kR\QÔ���M'�I�d [h�P�.��"����vz��6�!:S�Xi_�N��2Ӗ��G�����[k�����ݲ���RR)�s��?W�OHX��[hτ8e����4�����r�dUWH�U�0\(l��������F�%ÖsM�x~Zz�.3�����5��"�$�5���f�\�8w�}�a'GXXY�['��ݬ.��ṈT:�[~�I����jc�qC��n�L��,���> `���[F*�TKIiEF�]��>^~��φOL�h���D���������*�2�[��7��W�5�X�K����_�N����5�f��<� l���]4�'�F�I�g�$:�4�����xԘI��]ӚuM�Q��/�a������L����������E�Dfٞ�A���堠`k` �~Nj
����^�ee�$��5�D�z4�(*!R� ws��Hw�o��C:�fGT R���������5�X4�Р��#����Q��i�j�q֥�++,��]��/�={6������rM�U�x��XD) �����LN���:�8�$[WW�"�㍬>�X*f�v�q�T�@��n�ϟ���Y�����Pє&B�nX�}kVm���XE+Go������X���V�p�邺��*-"�?Zi���y�J��d��+�x2�%��Y���X9��c ��ڣΆ��<�@��7h���\dV���7�(bN��lh_�g3����J���G�B)����J%�~�x��������sjD��+��&�c�B�ވ�$8X�^W�Cwi{xp$�֑g��`(���AQKS'#�O��^��yTuG#Ͱ�s�"���p-M�E/_�����5��ε'�YB�x>��C���|c^v��z����?)�f�!�!�o�jo@�y�0�8�bicx��e��\� U֬d�)Փ��<�P�֪�Jߒg֘kۤ�I˦�JϾ��Q��m��Y^̗�w�����/O�Dc�[��,�na��:,�C��GS����[��o��Y�;M�^��±�*�:����;c)u1_o.�1��������QQ���%Ml��/��-TU*�~.�K{n�p��ȑ�B��.��Å����,Z�u��5�.L�nIz~�h}����f�SD�u-pu���XO���ڗ�(_����pA���L�C�]l����LU+�"l��������ѓA�_���	"��#���%��2�2Ӟ�JA�t{آ��),aT/W�,�������;��
V�b��RB����Tq�F�s��{�޺.������?e�)��b�������t!�D�1P΍�*?�r�(J�,���g�Z�=�����ɺU��F�~.�p%>�J���`o��Ʈ?E�¤%�!6�@Yg�"�jx��խ�G�f���Xg���}����Q�������	�2��J���S5���~���U�%2���^�����ʛ�hS t��*�ۖ:��*��ٓ�1m{_=�\[:"��bar-��NH�����ď���"���D�d����s&ǌ�y�t���v�66H	����c��h`�m�y|�~y��ܬ�oV('A��>=���"{���ykc�fD�Lji�A�o4�c\���kn�Tт�4���M���4xs��rx�4r�Sc���Hz���!� ��]��L�C�O�^W����b��㛥O)#��Q���9ؑ��Q&�ӓ��s�bģ/��e���"ɬ�'c��m�%�a���l��wpbS��K@�&��N�gD�)�w�k���V�z�/z2l8��R��W�M.�ķ�����'	���@Ȟ��8�a3{�9��ۋ�M��S[��-�WKǵ��y�5�_���P�Zk���VYi�*��W?1f���!��*m��3�q1*_�\;�ؒEg���X�:7�q���/
sH���9ѷ�\��6V\�p��Vʪʓ}����ˏ5�i�NIW]m>�� |��� 'N����sԃ*�$N�<�=b�;nkg��x��1�<UuY�X�V����oDӏ�dwť�pڃ?Q���Z��*�4NB��=��Qǘ��4�Tš��@���4�}��H%S�l� �l��lO&���њ��	��'~s���Ri�|���C�w�37�$�C���Td\yu�_��L����$3YGL��C���� �&g>�.�����)��&��0>�(�⸓���V����XM�+�+��0���5�&����Vg>y��o��*�[k	`�=��_����W�N�,����j��O��CT\�����Mwl�=�(���%��>��I��s&&�v�I rJ��U�e�k��hT��?�(��;���n��\���6[G4���z� I��礖[��4,�[�;������<��F�&Bi�.Gww��[~����0\!�fUŃ�7v�T>2���Y}�i��G�:�}��=�P F_bT�1��+��}]�i���,:�C��]b�����c�^�^lޑ�/�.������G���l;���4xm�6��yF6�܂1�}�@��-ik)�%/ƍ�#���O��S!\��썔\�H�Z�D�wG��/ֺ�>P����Ko��"��v����z�R�ԸH��D����%R fx�x��6ְ[,����ۢGC�xA\<���[�at@A|�EEͨ���_S�@����e2���l�ӯ����;�;>��C8\��5s3� �R�!���ܜ������_���w��}�:����SL8������Ot�D ݗS�
�^��Tϰ�2�w
�9]����T;��,P�Lc����,�BV�2����I�q�իW�o+&����b�4ClR��$�"�?G҉)�{�r��{Y�o��r�������IӘ��:�Y����Ԋ����
��1��R�@,�G �tCW����Q���)��9'�e��U��F�IQ��Mܳi�wnX��P�����T7�O��؊4{��x����qn{K�J�^��y�Å45Ӯ��:]U��Eg�@'��W�e'�l��2X�i���-杙��ۂ������9���[;N�u��}�:mM�E�"�>Tz� �����PD"���S?Z]��IN�W9E7��{nn���'U�
=�i>�J�
�����2�J�&�9�'� �J��a\o��O���y5m0�&� ��7���7JJ�p|���8P=V��^z"'��п���g�`�`%�(w���%��W�/*�",�rqQ�?��z&�ag ��ͅ��k�q)'��h�µ�f�5һ��K23��u��%[������|+�5p�{Q����7d232��v�v�/���[��)/��l�잸*�βQ��31�;�@J��\�@�5���ϬՏ�5L\]v�Y��ز�9�B ���Y��7�61���D����ۭs#(���
9��S�.���.�;@�D� ^����w��=ȱ�:$w��V������R�=���hص�Z����IY� �h7-!&-�(M�(-�(M�-��&�v�/*Pb�Ґ��C�1��^/'m��Њ{Yn9�d�����LD�R��R���/���w�%���1l��2]��'Mt9��k��n;I73�2� ��/����S�\f�x��_�]�M�������ȕ�"�l�$LS����{i��ɋ"�s�;���Ҳ��m���`0����2c�(�,� `��9���-Շ���������|�+{�ό,���9���N9$㞸t-�n�,�P]�zvv���W�	f�I���蓵��)����Ӵut
�?['�yb��hh ��5ͬMcS?����͎���K>z�S4���˞z�X���p�<�w]� ��5N���/���)�8z(��1��V�b�7YY�Q�B%��ea
�uɯ�`h�	�]�CT_��~�� ��U��Ҧ^F㫘
��h�$}��V�o���Y&����=<ܒBl�h�s������jk�^X}��C��_cA0Q�gK��{���iOZ�@���}��aɖ9�^\�p�Wc�P���QVV��	->[��(�|�gB�#����	�Og�����b7�ucгL�+�9��}�)�T<��uO�bN�sB��Xl�ᯒ��/o����1%�m!��
��;��[ȸ⧶�7]51�on=ۘ����,�Jc䳛Ӭ2����z�vR'6�34�;٘ +߂?5�h�K>n)�I���U�"�ۡ������<Hy$��]�?�b�*�V��/�Ԇ�G���4���#��/�đM���$x��x� 2+e)Dqc� `�j�� e� i��o����럞dm�g��Txm5�Y8C;�/��
�fs�Ԧ���N3]v����+�|V�К��s�<1��[W)�rv|ثG�ir��<1��~?��q���z ������'&��K�H��iӎ	tN�<���C�NJ����B�#���qx�l�:���W����Qvz��}��lE�~x7��@��d����T9�R'v��5�x�ڼ��1b��sҳ{���0�SA;��ʺ�Y���o9���0�W���ӷ���w��7�-滖{e��%&�� X��"�;���<���p�g�H�v�H?�->����.�o�ɾ��xG��RrTǫ�R��`K��8��u�YI�)F�9�ff���v��������q��,�ʴ�N�D��R�qW�y���>���r;������__H3����:V��4�ބ�~���6I�dO�-2$M�����RN��.���B�U����w����'ؓ�6���Q����zZx�w!vn�*����s4�v����fD]`���ä�s��%$o��zqf�?�o�`t�n��f�̅�5�U�.H����!=5!G�"6]g�"������o������^h�{z{~T��d�����T���l��3"�/����,�#�Wz:�Cf���+ր��k�1���/�n�,,�3*�s�ڗsm�--!���U�<R�EM��Yg3��Ɲ�Vwu�\/�#��/��B�trr�'dǮ�m�/�.R1�F�b�n^,������4�v�<����8�#��x���c-�d��k�4?\ln�Fk�q���|?��{���|�������P[�2�d�s�����Ǹ�_vu��`|%��`�b|IK9�>��`̵�k�*��TM��?.��XЇ��"���±O_T\+�c=�H:�N8���o�zSN�����\e&#�����.��(oc.C�-FT!�[k�D�Q�Cu� S�>M.6�/�Nj	*)�c�y+�fљ%)+�MW�bW�f'�'Q�S5H~0�	'm�j����=��[S������l�K���mOr��ƬV�nJ�vdA$ZH���@G���T=.k�F�K\�ƻ�d%}gV�MԖ���S:Cm5�
��n=�[��9�t�SNM�gнYgf��ga:d;B�;��%���b�=,:f��T��x��1i���/�LFE��_��~������?�}`����0 ��3�v���Ng_���ם�y�ʜ�dZ��cF�r��bP�@�����@�0��~0�g�c/���h�r�̌�t;V|�o�U�uq������A�v�zc�u�4%�P�!G#��gg��d֫��"Ͱ��g
!؉�li������+���60�k�3���gy����y��`����9|�C� z,-W���W���H�I/��`;��?:n=�3�e�h�1B��z���`NY{��6�9 *��d �`�֖� �Ǜ�h�ء_]�`vL��g)��SVL������3P�.��}
�ea�A��\�j����n��`��k�J.<m�	�6������Ϩ�؃����������'{i`�����өy����;��O��k���8�s�f��8��B�$`/[� �澜C��h��+\ݮ�y�N�Rp|�����xjwt+p���W8y��O]�S_����Qv^ǣă@���<�1sU���ypg?��Nޚ��$�6{���v�9�����u�F���xI��hifZ�]dpP�n���i�1�R��G=�:N[,���β�q�����a+绛kg���Lk����<w���<cc8[��;f��g�v�8Y�.,��(&*���j�5�!�D5J�l�_�~���﹟
㓀?.���3Łu+>L��=qJ�
Ӳ�޻�?e�QL�+��a-��әҢ烵Y���v}�4�`��F'J��K�S��*����8?O��.�������2k��̺P�D̔�P~qqZ�EUb�"�I-)^YzN9�[4�Wb(Ki¼i��}����=TVt
��b�0Q��,�?��hc��\85��c�J��M�*uވ��"��h����^����� ��#ƿ�߭��0yasA?4�"��y��Lp�1�t��|�M7@.������g��#�fL��ڴV�5��
&�/6����� ����9�՞),D��#`K~nq<��N�����=�Q��r��3�cH� ��v����f�E��0����3�e��<�nK�r���|CߤO��_)7^wI�j�T޷wޑfπ	,�9���VPP�@���]W0:QIOwBE5�t�ǯg�,��?�d������Ga�����8���������j6ݸ' !l�M�'V��J'(6z#;O i���δ���q�̀��j�P���R-g��b6)nҐ�KC(�e{Պ�7��������i���L�6K��y������)�g��f�����#'̵Fa��q��@���-�P�����a���q��ȇ���u����8�T(�f4�d�h����R�vܒ	�Ɓ'}}�v���lAR�F8K�D,���ރ EuN&�4�� ��72YN�ӳ��֜�e�)+��ĝ���l��7���1�)(�7��V�}����,jy�1{����TT˂����W3�-��9TT9��D
A憘!^c�Q]����2�`RI�����F�8�s���L��x�.��";Y�;O��X�Q����t��v���'�J3�b��ơG$�ZE ���p��E����ƫ
�pٝŦ�&�z��kٚ���{3�ן{�:��n�j0<8r��}R��K�n�4�P/�Z ��yx8�D6#����3��+d��T=d�G�2���^c����8�P�u�E l+A���z�Ų5}�C]��ʋ������C=��oő]�����2���\��xЉ�f����Mb>N��P�������e�C^�|��qB�I��StH�9_��\A:.�kR��&s��0��؀���Fk+��9"ɺ =Ҽȗ�h[iy�����je_i��l�����F{�+FH�*�9��^�iŬɎA+��$�h:x'��f++��U?�v���Ii��������I���Ur"/�r��zfM'�IM4%���e��jYҷ�e�7��q%O�Ctן���%.pCr��u��>�B�� &	�T�G��P�b�iv�����\A,�l�Ȩe�n���1o��}6�$��t8[�e����{Ϣ����Izr�\/2�"�3ѷ`�'����Zv�;{����7����W+��%	>��?7Lr�X�!V��g�.k����&Cfe�v��ۮMuK\�����Uq�������?���x�B�� a�?1�T�OL!�Uo?���MTU�lA��Y0�`)ջ��ie�o�!SV���kb�H)��Qs�D����ª���kzm�_z$+I#և��W"{����� �e<3��8z�(\�:FM����Q5fvr�����QK�tA׮ )��$�c'a㙾������B��������Ѱ���M&���{|L��I N*��n��Te��@��ʄ|\��rj�y�	��;�<�]�Q�1���ǽ��JpWۻW�$NĻ�.�,��hx��Ӑhb��HGJU�*�Kkp����g\���]8�I�"��������t����y�i�ػ�J�<��y�&�!�p�*+��BF�[a�v�xz�6���/i*��Tz_�f�307�����P'�V��63�ʳy��S�Oߓ��"����#���2���kpv�3<���3�:T�x�v�JџM/����A?À`�q#�E ��T���kjY�z������jI�t�*�>\d��
I ���o�3x��_]��B]j�-��УZͽ��ٹ���,�R���]�f�=?^�`���<���ߨ̓?e)��R�''����,��u�|���
f��.;�}�_���J�VQ
��yrFT� T���͗�X_<ͶQ�oRà*���W*�w������x
�s�&��	g�M��t����;7�!�R�g1c��n����M�F�����׾&N }r���@��i
�Z�x��N{C�'1`���Ϧ�95��Hym��<p�ј��5�/>�l�R�0�3c�)ݨ�Ȍ�<�� �`�����4 nIea�?�1`VEX�ɴKL�b=�]���t{RԴ�=�r�7��V��/�#��a�?���c�`4�����ܽ8ͦ-̶U_iS��2�&�geLo�n�g��Ee�����9�0�J�&�'B{��=y���Zf
��2q@T[�Z���lR�j���;�k�ǻ�dߗ|#s)�f���ꆪ���O'�m~��Ɠ��.k�jO�)�:��������k
�P�'�G�<V�ÿ� g���y��S��SN-SK��-�@��uD�W���5Ͷ�?��FW�r�Z��� A��c�6��H�T��Mʯ�D��a������͸���)��IQv�EH�ՙ�TpZv�����[�!��7�)O��
O��ʯ��x��u־�T���`���o&����������]�b�ȵ,V��Afw�o�!�⾮W��.]�
�aQ}���(S�EQ��) 5 � �����B�մ���

��?F;�:)y�Z�֮I�Ƽ{����&�X��ĩ� 7>�Y"�k���9L |�c�	ƣ	&�)�Ƞn�������6���n�Ɇ� ��ȴy�X��V�@�Gk5�)�L�¦7ަM}�c^�b�K�4�m��)�[���B�z�TG�Z�о65-�01�����Hi&��h�a�iB��G������Ezp98r����/9t��VL�U��������*D�Дb�9��7��=��69D�g��_��)�̀-��:n�!I���B�Cj<�p���s0#��9�.
��/7�L�}��Q�M�*�G�c1�]&(�_'*����-��{NV�o�@i�QyPN��o$��ef15����ӫ�M�k�
����s�Kmg��L����!S�4����"%�ͧ$!,I�
�I����Db�ru��=���g�w@z^0]�� J����>�c�B�+�e>?ʯqFw���[�ϖ��fژ=�� >-�G��S�W��oɓ&����K�`�NX�N���zRP���9�c�J���\���>R���;-Ast����wx('��Y�;��v��}�0A�s�ӎ=�r�FJ�S1�QO�br(<�S1��ӤR3����X�[��F�[�H�X��7�r'���n��`��.iSL���r
3%���w����	u!C��m��ÿ(4������pz��0u���gJ�F����R*�M��M�x��yk�j
q�݊��h�Ĩ�qV�����^�?Z�>��5��":��,I�2�۫�w�ϾT��A'�)H <X@�%���l/۴a,�h"l�VUt�ٰ�c:�j���5�~攐�����8>��[���V���	9�W��_C�x}lz�Z�8� /��o�U5����"���j�*��	��9�����6�j3�u���UC�mZ�B�3�?�V�9�=FwH�sڋ	��`Z]����ȣ��ڱ<�lt����i_OO+��"uo!��.��Ƀm� �K8#k��f;�{s�|j}pl�sX�JOM@��v}�
7�2�������K��c�[5�)�򌧜�]�������S!~�Ie����#8�p�sUaLLL;XY�n�x�0dYC��
uo����;T�d�m��l���k3�CL�5�����Z)���.�o�k� �T/����m���2���o��]�UqUa��T(��{.KAUV�<h)�l��E9�R�{L�:O~x����A��Y���,z�Q��[As,���O�o�
1�Ƕr���W����v�>pq>���I^���uLP�}��ѵ��������[��_��|b<9�Ҹ~bSyB����t��VF�`������,��T`���r�.��igx�4I�}�SA"���$�rg�� ��yUL����7�v�M� �����S��ՅŮ��%�D��Vc7�nKS�l:�jLCD��p�t�
�hpX�J~��Ì��C����<oG���u��A��/j��'
*|��L�E�.F�JA6��f�*�.FG�~=KA����M-�L�{�h�}��/�y'��� w��|N~ /�+ϱ��	�vn�M��	��9W��mzӴR;�U�Pf�lLJf��n���H�IT�f��0c�bBb��>f)�kS�c���,�w.�U��	9�B�:�>Z��w#̀@���b�q�E�M�J]�c��l��gչ߻�[��t�xٌx�{�M<�UK(т��1���8�2��G�$�:�Zd��Iz��T�������,�#��U*+=���)�j(���]�LH�o9�0�̰��Վb���� ��A|��A��}l�*�V@ ~w-[,��tFִ?3���U�lz�����:��:������R����$����D>���zN6A]�
�^�QIЇ(Ed�Y�aRS�i���7u�ƙ�5\\Bb��?kve<�Ol#�X&�10հ���@!{�=A߬����}>�m!��H�y8}�<�G�a���	-���熛I�^�1M�-)h��-�3�-��g�5�5�O|I#)w;l�� ��?u<��,��~Ӛno��E��]���� n�g�#�WI��������Ku�
���\Ӂ��I��i�P$I��뤠��;@,���8-ױ��iJ�v�Y..n?�:��?6lo�4�e\�=�hͭӾk�'�&JU�����6����!/�q��p���,�NG)"�<��h��������#�����jfh��Jf�l*�[!|A��� �*�wS&��>����I�x���tg���f�k��w�[h !��:��O�^�9-�$7J6�O��v�E}�Bd��hB/ƇormR�F�&9�G�<c:�ri�3p}/f�4#�� i�*j]��YX}CC�Dٳ찲L�����Z ��ʽ��Z>o}�Z���orr�i�!i��\��ߘNмD������+-�: v/�m�H��!A� �X:�{�]{QF��BO���-�u����'�U����7�RVF�PC<�o��k� ��ş����Wk���D%V�2�{ Bd�I\s��R�F(�Ó[��� ����7�L�}�nq�y<|�i(�W�i��������g\�����b�+��>u�����苫r̓{�ȵp��&��� [^f��S����:��$2��F3�r攺�����}7�R��1�G�����y���������je���a��#�8(M[dv>��s���*���1���ǘ�vw�z�L��ti	�x4*�[XNc�u3�M�h�Q�f����	��;���%�o�g+Emi��H��|���J��H��p���M8���a�G�k�C�G!
�����������~���Ht{P#����V�|F���䯑�R�|��[&����%�Y�;	6��@+X	LI�� �_�c� ��j�q�qFKrP��_���g��Y�������/M�ca'K}�����u|��u63������ݯҋ����^o~v�"{p��w�ɞ`b�$���	��Y�lyt�L�Y�d=[z#]X0"�>�S(;n���a+Ol˪��=oAp?an���Wt�+���q=�b;�Э���TT8KI���Ǳ@���3v�qU�)4��o��n�c� ;��-�\�j�\��D�8}<��d_ܴEURP��\JW{�4���U��=�9_2�RK�@���������j�����ɦ���,=m#�����m��Q �3�w5�o����<q�R����Y�.�L����*v,�����h%R�a���6����Z�E7#X�mZ���.��p��Ն<�4�ns��N�!�0�M�`Z��0^�0���M�r� Q��n�������������ox��D��R�z�B��l�'�z�8�.��ND���z`{[�hoYd��
�1�=���/��:���M��R����(
��BM�D�$�%�d�5M�B�ވ�gYBeI�d�ٲ���;������3�y{�^�ܳ<��{_��)�y*B�f���K��������F�l���IIIFj�ed��߱��ח����Htkcr���X�^=�e��.|��� ϐ��e�ofX��Lz+��x�s�b݂gF�%��;<�ڵ��*׮��H���PMM�!��(J��Wod����0����o��&k�^9�?���Pc0��{<�\g�,��W��}�Ҫy�c��j�ո	�lƑZ]�u��n��Ƙҋ������>>uib�1���� |���h.ޯ���y�V�鄔#�I��r�u�᳻4D�t�T]k3;���������Θ1���v���ҥ|k������Y���u鴤۠4n���b���%����}�z�#՚����B���� [�/u�.&&&Fmd��}nӍ�T��d�l�k��4>Z�޲�%:�bb^$'>s�v~����������T�.��/�n���ԥkH�~�������d�	6�#_i-j�di�L�~���9�PR���࣫C-�&3�dŗ��Ō����Y��1���.���\�LS?�k��K٩<�N��h��z�7�Y�h��o��M\j|m"��%7��vJğ���y��Y�ً�n�)2�;��������"^7�:������g<�F�q�)~���p&�"��'�Z\��<g�6��1�l�����J9S�n�����W6�j�Ƣ�j4�_87X�LD+���tkLOO4ۅ0��y=�Z��s���t:`�m:��t||���=I�Ul���.�����_��s����ӓ�����o���ï��ދ���w0G@�.���{L��q���W�D(��=�s���/���=���];~6��N��/w��U,�n�j�d`⯕��.�Q���r�{zD�����9Y�-vx��z6 �%~aҚ��9��RJ�� _0��|+��c��]Z1#�w����5L�Xv=zd���B���k��,�v�P�Ն���v��5�w,;l7����*7#������q�y[���=����[��ol��X�����F!�4���*�OT�;����2��ܻـɩ*ߎ~�H}ˋ�]�@\J�<��·� Y��J��wzys�ߟ�ΎU�d�<rƦ�V|��]�j���dq��i�l���u#:�����M�ͫVX�V��Nc��_�����*/`��}Q~#X}��3Y��f�l n�����w]^4�o,;�`�_��6)8�:����@�L]uL�^���/Y0�J�~����y�o�bzƇ\/>��� ����=Lo��!.�=&�-�����+拄{��Wy���H�o^�`�ӿw�8~�g���6�:���/���Zt�*>�\����*�\���:rݰe�|����c�E2�j�.	H������ᙙ�/�}g�9�M�/�t��L��,�En�2���;�&!�c�3m��@�v�O��y�s\�t2�o�a�K�2no��-g~u>RNf^�������m��y~hP��������
5^�������%���/�S�%�r��mL28��-�_S�-}`5���l��\��sms���#w,��V�[V&B��Kt�Z'd�c��@QF�Pѡ���?d:�?R���Qxd>O,+��k�[L��x�8���,y�n,�h�i�!����~�����ꐐ�f�a9�n�yќ���,K6Ez���ױ[ ���
�\�xHm�Ȼ%�

���q���vC-�w�`�9�������(��)�k�~�L��|c�{g����?�׌��Ͳ�O�j/�tx�����=T�	����F-ZC�9ӆ�>���Ek��ۜ3���-�r��\߇aןM��\G��au�G�-�7��	d�ճ�ۏ#ڿ�i`zd��ЏG�wx��άʙ�'& 	��#�k=�dr<ȱܠL[�*=ykD�,�@҈۬�����~Y)W����.r�,�낶�t��8;���ZɆ�S��^[!7�'��?7ƒ��a�V�.�g����������ٺ�+mQ�v?�8�{�;��}�ï����*�X����W+3�W�i�l`z�L�S�%wy���������7:\F�rOrΙ�Y�cY]�A��%�IF3�2�i���<#/h���������Zﶁ<.�o�s�jD���SAY1;��s��f&�����"8 �&�*�8�rGw���Rg��m>=���]�-�-O]�9�x�i�SwG��ɱ��(h��p��Z��%�xf�~Y����_ڜ�·�bW|��?�<=)��]�Z[��M�,�"�BdɫrEO��aW�>�c�� ���Y�_�.��:J>��z�
g�9����tk|�my`|���\c����-��ba�M
W(ᱶr�cꔹ�7���S4��*� ��E�N1ky������O��>������0�^S��yӛ�Lҋ"_@�zmj��D����j���_[�V&���}}�.ݬ e�쥜����?��h$.��8��*���:A��;G�\�g���K1��*�U�w�o��f,~����Cf�92�-o��;�q��R���(��e{�E#�k��*�ҕN*]��t���9���,��x���&<=/O���f�]��,;�t�jHB��G��4�>m��O��"���HZ�,�]�Ƚ���v<�5##���Tt	�e�6;5^g��\��r���x���M,9�ԝ?1�w���B��H���RR܍��Xa��8�����������{m�m}`xFZ�G]�u��,�Vqu�20)�a��fYܛ��^��,���h��{F���6(���Q��rؙgZ���DH̓C�a�]�R�t˽��Ѿ߮�վ�O��E=�y�2��1���1*��:�#%�����6E=1(�$���~��ik��3�|�@� ZO��/�[�9����չ��rS)cm�J��M������i	�1j���"����of����
���14-�Ѽ����8v&?Sݚ�n�%<�\%X:@�r��X�%K ��m~Y���q�wtW����d�/p	K�i�c�4~JX]�>(d�ޝ�5�~W(L3���9�X�dĉ-��ϲ-��:9'u��p?X���Af�
I�'I�'ܷ}��(��`Luy� ��d��a���.���~4[���aE<|������I�vF�L6�:K�9��'�@�G����/8?�d��V�&S�Y��,	K��@#�4�0'��k���u�lw�	�[��}ť.s��GF�x!��S)t	;SL�V����)3�i���g���OoD�/hL'�F�p�xk~�A̯zg"����z��3*Jp
}z)��Ѣp4|�ڋK�w��S��1؜E�����`j0k��$scQ���@i�S� [y�s�1����5Y��|����(��H@����J����g�r���鐇`�bo�Q��5G���p^c�(����h� 7!�E�022�oL�����S�?5�S½�k|���i��`	��;._Xf�WVZ����+��GWY��6�B��ɓ�z������i�o����x�8�/ϼ9�}zbH����г��@�x�1Hr*2/���O��he�X�$�� �ffJ�'����h-�(���VE_���"��^É�1#S�*����>���6Z�:�.�,gn�o�g�u�(�Ýa<x���d'��lAJa:?���%���j���_ @�+�z���'�W���gn��N�(v��$��i�O��W��9���Uֱ��׵�LRz�L�SR�����u	T�-�5�w���I-�9SLФ&��l��`��_rI�4��+K�y:w����K�kρ`\i����P���p�f۹k��:��i3���"��[���W\��H$�3^Rv�Ȗ�"����&[���V��n5�
����P����m�	f,a݈!sƟ'�`���Igf<���$�"(���{m���7���[�(�4��_�c�Hd2rt��j���6����S;� ��D�H���G�=8!�+�!���)֜��Wn���J�cĥ�<���̕��x�^UUq�^� xD��cl�����r��>�����[�)�;Z�}�m5l��x��]�:\m����|���z���H8�OE��������O��n	�~m���	r7�E��5�>&Wc�L���JR�n��rc�W���u��6�/6��С��ڨ�3�;@���#��2Ĉ�A�J�I�ٶ�6���aT�UU#����r�>�sދ�	��vt�~UQ�v�A��?���Ul�qLi��6h��[�Hv('���%�_A%	��Vy�:!��[� qT��ы�E��8�%XE8 �E�;���Ȅ�Waҿδ��;��cvf&�_�H����K����;R���V�6y�NOѵ�Zl��{�Nl@��u"ٸ��U��샲;��o��hGx7NRU��V�P�HB�]��Q��Z/��Rp��Ԏ���{r�W��㾭���Ub�B&���H�!�����_��Fw���t��!��l�)�+�rg��R�����)ہ<</�p�ۅ���o��*�L_t<���"nU���#I���w��� �(� l�����@_�~Y�y����Zp���Lk�S��Q]>���=�8��~�צ�U��ik{@&:��x�h��'�����=Z.E!�~Հ��3�[	��x� �$��0��e{����P��ޏ��'�g�5R{΢��V����8�
�=0�E�:u��X{$Q�b�^���S�!a�t���n9�k��s8�NP��lB�p"�3� 8�̔�llB��B�h_'��IZ�+�dZ�a�NB���-��h��.nt����{�����"�:�Y%�8���0�]`�/���5������{�?��)W��g�h�b�ȕ���@�h���p�u� qm�W�Q�b���;�	&�?��J1�P�+5�YMU���5���OJ�m��Tay���������m��<M{oJ^?��$��t�%�@:ݛ.eG�|u�CT[8T-��9������<�.���T~tو�3Me��:�8��G���i��`����w�m��٠�>A_����R	W���&8��Q�eM�� ��γ�u����U@9��u�ƛ_�hf�*#�����h<�	@%�*!7��-�d=������T��?�Q�6����n��qzfB\��W��D�N��"�}ޱT$���s����bBP�UK �����.35�`�dީr��w��h2����EP�?�_ߘ�W!�,�5!B9l�ξ둹��E��9�9_z�l��@}���y�C*3��Ӆ�ڇ�/�L��#]����[�NAݺڢr�=�����7�;��`��Rs=;�H�4� k�z�E�U���x&a�G4�j{~�5�==���J��?	�����q�P��\ߦs~��v�C�&%&�'�~n�*�C��S*k��uN�[iЊ���AO4����H7`cERCُ��It����o���j�����q��\��G��FiA�
��p��({�0�l�ך��@�d9�j�
fH���]b�l˥48�;�]Q�u�ŏjG�ȷ�ŏ,;?�$|湚?�y)�A� �|P���"_�7�Wy��W�@{�[1=7=���+�B_�k�l/ ��Ϳ�*<uҪ�#}��Z����R�x)��E�yL,�Dx��g #(V��h�������T����6XHc�~�S��	@j�:,���/J����E?;Ĝ��;>}S�:ؔ��+�
F��rJ��S����k�i�����m�W�_��lGF1]����o	�.eR��">�������]���� y}H�
Ņt��wKx���{�Hl��Z^�K�I�S��i����*�L��@�5�ހcV.8�&>���E���;���ہ ���*T5�	�-z�`l���Q\N�7�n�Lz�����@����,L��Y]�:M_��2�y&�b�a�b�ؤ*7��${6��X!�^��\�H�����"\+:���m��f�n�sl�L]��F�� 1-?֋��xl7A���ȳi����J^5�� ����$��U$C?�r�w�oL" ��Vޑ�C�m�Q���t��_���`��YH�AM���H['ʥ��lX&��x���Rrc�|��@�Q�m�j_I��أY���B�= ��+�w����7����e��}}�~U���F���4���l�4�@z,̰�g����H�17�R�_��U�Y],�9k�Fi���JΎ(�^����#\뎊�B&U*@�M��O��[��̄#�*|����ͱ�1f)$�}8K�J��U~�5¡1�o��^���;��;�@����_r36��ƬAA��l�e�2,1�K	2���C�%LuY�7Z� �]J(��d%ˑ�PRV���}5>�"dJ��"<#H����WD����b�W�M�&vkm�g�+�L�2�T-;��5q&���N��D3��vg�T����aP����bc���0_oU�cD��j��D�qe�v�N�2���n��/���V3�HG�����f]�v虜�,2R�g�!�'@KE/�?Z�B ،�<�&�ylT�i�t9�=�it�cEe�(�ȭ�$ mF��졄P�[5�gF�a'�Z�q��Y�ϳ�5�o_��ӥ0}�Ɂ\�1��, Zb� �dL������*�4drCqZ��w�[?"�����.���j��'ٔ�h4�����Gp�ȳ��[t���'>�g�����魮A�L����x��=�҂�1z�ǳ��{7�� T�,D$md;/2?�]��w�ژ9D�����觗��l�gtt�x������-�>'((�$���n$�ð�"�(�]���{��0߻ʂ������[�g6e���ת��&T��Q��`�8�[e	�%,�+��񾺎�hu����Hv/qP�£�|�
�C�M%��[��.���^6������Ծ������QA�!8`���?P�ʑҲ��y�Unʙ6/-/�(w��$K��G3�٨���w�v��I̔MV$ e�0�H'%�L��s!�$���%ؓP"MsZ�^�ƨ�\�G��1�"���R��BUI�V����XO%��r!�4�lݿ	'L�����_���/���d%<ܞo=8�y�+���D���񮝩�+L������Q�ǳ7��`���v{�`S�x8K����I��@��4@�r�k*�D>��|KX�fV]p?���6(� V�T�w��M�CI&� �Yv�-�,����i�.�<XS+�Q�* j�D�8�G6[�����L�"~�pZ�`f��{RSf�+N|`Ү�W߀O�(�%)k��[ۃg�6�\gF�@/B��̞n�,!|�6�����%ȱ?���Q[k���i�T���������>����� Ly�X����"�^��R���k\{ .���� ɝ4�B��&>���}⸼�/4v�DF�����QZ�5`�r�� �#�;e,�� 
��'jD֗�O��Db���*X!{�hL��bv��X�RŹB~�B��2?񐔼-1O�'Yf�B{������0�;g0q���wl`r��D��;�l?�b���Ͷ�����,vV��9��\<��r��-��R��د�qߩP��j���O���>�/�1�,Ј�M�&� )�)�ǧ���ԏ��4���j���h,P�O;�X�wy	Pu$Yu��ʿ�Q����=;F��WWO\O��y?���v�$ڦ:226V7��F�Ȁ�l7�fLd"�r�H�ҽw���m���-�6���{ ,��jv$1\�FZ���
`��Ϳ�sIX	*�8��s�˖�N0��ig�D�ς����\MT ]�nÚ�x��v�anO�����ݿ�x�>�T�X1�@��'\_2��\tצ-���Hd���h����喽_^��Lu�����͚���0\J��~�9���7��&�:g��S���3fgj|�fNA�]/��q��{�'lv,t*V&X���߿�hI�w�_��la�U�����#��6��${�f4�&dZZ	�'`�N����1l�����"�J��!E�|�5��FFۑ��'�`ɀ��Z���4jPfo����]�g����������b�5��B��5b����[R'GM�x���R����&�0�x.���h¼U�?K��^�>�E��އHzh�#_�Ep}��p�6�}�S��I�N���߭�&�������8�L��uI�a�5M��~5��9.$W�w�-�Z�t�(���4P��·���' #mu~� ��s�]�$/.Kފ���W��qS������Y1�!�8��W�v�z׀j.y�y��W�g� �n�i��Ͳ���V�x��=3{�G�ǰEZ��0��l0�jȰ2�Նr��2R_=R��������@c���f���ysm3*;�w�災%�on��*\nPF�^��]��O�" S!#��8�h���:w�bx�
i�_��]N��	��/yksrb�%�	����q��
~{Q����Q���ݐAmX�a��?~v�`�L��wF Q�}��A£���;��g��6��A�Y%��e�p�Q����k;�$a0ʢ:01��`}���b�ױ��Ó��~��@���K�$Vs���>8X��M�X�&ڋ�LOx��ȝ�O%3c�}�-��I@�S�bWFt"(�e{o"������LKpYٟt�X��T��ǋ�~�[�ل|����+����3����U��"����>V��G�K6�)H��h�q#��8���l��ɩ���*�}:�l�dD[v~f�hm�au�{�vG7���dS�b�׷N���k�P�xı��r�tjD���>��G@���˷B�^��2�F�Ǔx����+����� 7�7V�٫f�y�@�h��/!�8�;Q�}��?/�X&�6���>߬��Q�#h{���>�wWߊ7a��ގ�rTL�@@}`����4Ǔ��I��:v�=�n^@*K��*!`̸���+xӪ����b\�M��	���x�>rc����F �#E�6:	vg��DLKV* ����+:W��vI!ԏ��kWi�o9�C0<���{��BB;o�:��O&C��9�홹|��k���զ7�3��b�V4g�	�v0�(�j��OQ�ݡt�+1t3��$D����h���� ��8��)�tVhcϥK�?ho���≶nUU�p"�F��k,	+q�n�z��:��{���mb���5�f����q�Ӡ��h���������Z�����,�h��%#���l���!_/p~_b��j}�Q9ܮ����s���)�� �u����י�rX���)�����ҟ�?J�Y��0)����<3理u�I�^ml���y��^��n���'ˎ�6�3��8=��P	_�f�XrR0��$�}"%k1��42ĕ�n�	w��dA]�Jc�_�P*��3�� x����'G�8�x
�}rrC����Vt%e�
a8�r�i7�`��+�-Y��(©49:�gK�ݐ�,Xn�8���R^&�lQ��.c�<�7l�28�6�C�O���| 4
��������;��
������4)��:DM6�n��z)�A>� �#bv:��ΚQA���eE�!ޗ�AK��$�����i��B����eSު��''>����e�Lj%�?�A���:���Ew��/���Q���]����� �<rɖ&�& x��ߚ���b�;����Xa��ܛ%
sB=�,:���ju|� ��Y7�:��-�9\��#�2Y�J�o�@��$kT�����������y���7�$~�jH���&��F4�_v%`����I��`JFת��T-�਄�9I҅����!��'�m���ī�)(y4@��pV��vk����/U.��;��7��-L�s������p���C�E�W��Ԑ|��F��QDF���"�����H"�w؛�M���Xh��Q�/�?���e�t��8�F,h�����"7c2��"Kִɡ@=;����� ���@��t�4�mw=�r��1�V���d\���c$��L���dg	p��_?Y1,s4w��7ٍ�\���g�Bo�-5c�nr��΃(��i�fɺ��WTdj;��L���*����ȳ�+�3	&d�SOȷb��4�}B�j!;�]ƨd���e�,�y�2Nd3S��.�9��_�:�ʖcg�-�W�{�#6�3!6���ur3Çѷ��y���FJ�`͗k+�i��z�x(9��qW72V�n.J�}�1�#�&������g����1�p��
�i��H��¡\~ҵ'^S9#/�Ӝܯ�8���Oӿ���ʳ0w�Tl���Ti���������w-�¼����MR*w��H���y��Po���V�&�^�kK!��j�h��-���&�^��N����k��[g�E���sPb)��,�!^���A�O%������g)������!%�󀾴�����VPk�?_���I֖˹m,))i�>��,�טq״I����;���+�-U�;�OC=�t���|�O�z,�Aޓ�3�$�_��kW���S�]f��?�Ĉ�(൏�����8�\��bdo4vC��H��f���7��gR��o���7$�O��T�S��9��!�!H�ɯ��~����v�7}��p�͙V�*3@�`���8CJW$���oN��m��r�{�*����ߓ���P��<�h�� ���N"o;΅h�{�9��477�
��O���H�N�A��oM��2�ID=���/L�������`@vٮ|g"z���ޚ�wDfw��;V^��8��< �q���@���X��ޞ�����󘗒c�~_D>0b ʕ��P�O"55��q�(=nj Ge�v1��t"�Y���TV~�y	����
��X����vv)0�H��.!�Y��[�J��ّ�o޸ͻ�m��W���226
��J
`L��H-?2�-��� �$�n�F���?6��{��ڜcֿ���ݫ"��k�Y��ח���c��">�o.a�74܆����G�*^���FI�: ���I� ���)�%*z����[�zb��yLv��q)�.��sr�ڣ����D�u]��\���� ��<J齜�U���V���hs[f}�S[[[�{f�J �"�,.Xs��tP\e��5R��^7���"bsy��%��.bN��"pd��hV�����;��d����\܀�v���d4A��\�J���߂�JC�#êƜ��j��o��CKpA��I�(�����a� �u�z�߮�R$���2�,���U��oP�%8��(�.�@n(?�_lS�B6r2d����J|@?X�g�y���!:E5I/�� c��U���^5fFĻY{e���'��?7Jۯ�r�
���+�PA$��B1G�t�Z��=/�S�m/���{����jO��%��M���9�v����7�V��N[�����f�I፲�ļ�dS�ɕ+��������G��bY�njnQa��i.�B78�����O���24���8 !VSB����Q&����?���^ݭ���������G�mNڼ9�<@q&$|A�J���mYK3.���TRo�A�{Kwi�4���˕��mETVH5pV7UE�v�ӥ�¤P���T��\�Uf��nl4E��'�,��B�e�wY��L^B�f�P��+�}�w����iR4��^^�輯��<�|�B��.X�a��`sI����D��Ŭ �$���5�q�N���0�)����ɒs�yO9lώ�S���h���Yy9Pk��~qq43�n�a9Dd��?L���.3C.���ޅ^E������/���b:�ҰD�&��������骷O{�(�w���r��9�N?�}��UܫI̲� �
$8�S���`�KēiNc#��gW�~l̲ѿ��H%����)����V�U3��?����7_��M�HT��7ֽ��h��W�:��~�|-���w+.:�N��O<5�%�<�j�'(p��`�/�����,�q2Z�8S�,$u������ �I��ԯ6 �#�#�EV7{����o(=ۀvI�u�O���q� Xs�~Ă����MDN3�Ej�Z7]	b����`�����$H:�.�m�?!qC�LU�[��H��MQ˿#�nZ����'ݎ��+���e������u��7�W
�"��W-,�L򐘄]SK��ۇ;��:Y`锛F노�k���v��n���	b���ݗ����S�6x�V����O$���ĸ���W/���7,_��yq����TF��TK���M5�����R!{�x������i�O&�𦬉��㛳��E����������?-���D�����q�m˺p	`�.I�ɑ����4���O�$��o~�y	��9r���N��`5^��Ϳ�#ֿBk������G<d�dj����$�;*�M������	o��^��sϼ��-č�m�ߌxn �� }�4��l����&E�ͥ塷k���E~)ѮTE��/��F�'�m���PT���l�m=��WC?T�Q�ڞ�C�h�m)p;|�`\t�T�����aH�# l�"�%cA�w��N��K��r�|[@����Y�C:��f�L����$y��6�^.o2��JUZx�S{�����C%TU'��&�+G!��VS&MPoZ��� 
�4�{���W�w���j�i%)�m�#�����ߜ��ͣ����>��i�K{B~ۆ G�� ���`'��*�&��'��z��ojྸ��K$=�d����V�5YY@��5 |�=4L6pPI��Iqߍ2^0̮�˨��F�],�k���	U2����WJ���`�ɂA9Ř��jr�P�y]'7��wHu��^R"5��8�ZJAW.�2#��ܣ��>]����RO�-r�|���פ^L��cCN,qj�A��7200 �ٵG岓i��Q�e���l�55�G��t8��&�T,D�?!�FF��6�;�&�#�� ���*�B� B= P0 �()R���H:ե�Y��oA�bV���Ѐ��/��h*�5y-"�qy���f�������*��w�+�=�a�v33�|�7�8�bU?��n� o	�~p�V�y�\d���/8����V��g��8�R2�
��W��*5�u"�e%yCs�!�-���F'\��{�W��=�Ž��o^�jr�.��`�uC<O�wc��:(���$��W���U��9�J�#��i�Zd\g$6�8f����R "�n}�p�.Pq�BR3�B"�Xl!d%�U�[�~O��_��Dk�Ϟ�*��s�X5�Z���8Gf����UBos)�Y}``���h�w�С'�b�E.a�L�d*ں�����_7��}��K����m�l/o�$�
��!���_��˯��R��>e�{��Y�nK9���P�n���n0��0�5!��7��撥�GX�h��t痜���ז@�rO� ��ᷚ"*'��[:2�!�u�y�))�!�(�=��Bj���s�.���k+q�k���� W��D�B9ڏ��O{�G��'����ɇ�6�?�����_d� �&���wE���,)�s9(X�PbU���dvR��˹�R7���w����0@7p[�ՕS1��:IW�e���L���_�P��迅��%O � �Y��P7I`0��7��C��'�.L��� ��Y�����ߠAю�u~�e�m��M$�]���V+�{L��1�o��M�/���������I��J ��з��wp��G�ӟN��i+�c)��C1�����?
��.���n)Sb36ұ EYL�^�7��u���?}:Ff���������ƌ�wEՙ�'�Bĵ�dv�Q����0���CAU���V:뭔-�L1}��su����7�����#��d�RX��a���^���u�A�~���n�Ŀ�`�6T�C`����#����`�r"23�M
?4!�=�O�p�dē"�e+�z��'kNZҕ������m�Ů�O�\� �i#�%��J��M�_����ad/�/������,*>�$���
�-n]@�klj����o���?�n���<���c�k^����}��������{�D�/��>���0�0�<��Ҵ��<�Y`z�+*�=9���nAA��p�7-+)<�>����ĸ"�L�K_5��Q.�@��vu���+5�g���o�e��i�#e���L ����V��|� �F��Q?.��4G/IH����J�%`&ޕ�����'�%��3)���t1/��4������ȇݿJ���T?��+܅�#��Z-A��3��q		H��G�,���!�\���ᦅGA��t|w��Ne6�E�#�S�z��lFvxz�rH!R,b�n�J�H�hf7]�i��d�zۡ�1")�֟��F��`R��X-��Q�W�^i�96��<�Y:1{B�p�`�_��@ 봵�?� 2����sӹ�R��F���y�/"Т'����s��HGQRNN0z�eZL��'�����P�����wzI%�Ԭ_C����)��g�|A�ս,�p�	�|>إ����>5��6�ih�i�ȍ�Nb���n��.痳�hnn�m٤�IMJMe�|����&�O������(ĸ���V�K��<}0�h_�sG�z��Y���;�|\\d�u��;@&,W<ȢY��m��#�����9O ����C�����(=��j!*7o*荎gڔ�e�1=D�����^��[�O��-]�M�s�&TKa�[�w�$����7cy��2�A�ڙ֯4����u���~'�`�����7D@=��Ө�t0� ����P���Sdg?�d�02�H:��

�r�����rvW� �ǜ��APxT ��N0�a�y���HQM�Yvdڷ�����.W��ICCܖ�fm*�RK5��4�H��漉0b\��P.�l�/�g�� _ so�~͵��2���h!(��X|��$f٧������һ�ZSSC �"�j��>k���E��Dz�5t�K�8���z�!9i��+W};��Y���L^�3.�K��X�*��z����dɞ�lK����2�s�W���ՠ� �ǅ�Ї��%��Y��B����aoQsy�P��c������E`����|X��S�fޅ�]SM:�n�QϾ�� Ϯ*a<��H-����������@����,�i��v1{��Z��&���������OB�%V
�:�������8�i�Y��e��`J_��|��[v���|�P;��ʧ�Y��O�.��jS��UVH��]�1<p$�g�QdA�7$n|xq����}T�o5�����"	�?57���'��k��Z�B��Zʵ��"UI��|)~�Cސ�2ˢ;�=��ב����*��r8�3�s�,Al��2��$xv��-�YK�6/)!| n;y;���`SF���!y�3蹞�����FQ�o�P�Z$%'?D��c���p�#�|�[�,�i8��,�Z��C��]x0{��؛���'����8��3�2�!*+�V�H�
�wu�.��!T��A���Ch:_�|������7�C�v�X4����)o�p�ᶃ���k�"#)M�HH�2���"�V	�1��!����q��:(x��z�|k�͟�S}	���&��"�z�1p���������B�
�q%�/&������}���t?�	�v9]�Q�|7���F6���@A5Nn�O�D�_^|���}�z����+��GG;|� r/ bYA}�t���d�������>�k���B��L�������/�k-_w{I�b���l=�nC
�i��h8�VVE_䗺��qj��U��'|�ȑD���ux��XB���) �]�%��Q'�h߃"�ׅ��F��H<y!�vI��j����M����A.y�g�ΛU�s�A�[j�"O��Q��b�Ή�2���i��°�u��KTBߗ����B�?����Oɸo�Ƚ�����*�]15&�I�za���p��@\U������#�WY)U9VC*�M�!=���W0UF�Dxu}]
���C�\ޭ7ZJ��[��xIÆ@l"A�*k�B�c��M|FRe=be�&��Jo��'��J^J1���9S>�* u��X�+$}����9���J&7;�}<�����Ѳ��//��#���V��m�=ڍ ���\�eQz�c [x��~kaCe)E���j�ܢR�jx1��9�Gn�o���n�!�p��?�B�W,���D�j��o4��8�]=�?_��p��,�̄�D�dxbL�}��� r�%r7rBFi���2�YP�4\��%++x�3�b�o�k�vus�H�#���B�x�1���	YY��eDR*܉���w���:�_hΰ�GL�K:72!������o��7�4E��]�/N~�8�� ��.�_�?��z�1E�)Ù�_��{dg����ri��[%LŽ$��P�a�afH@�����X�s��"7<-y"T�����J��a6⸡��۬u,�C�A������#���O�<!))k���a�4�-0�L��T^�F$���"I��t��n��C�C��1 ��>{���|+^�Hm���,�@��Һ�V��z��߆v8<��Saɢ ��̃3*g��Y��@"l�Fi����𸝧,nuSs��G�e�I���`�,�Q���A����!����[(A�ȕX��H��Wx�Ȋ'!Qkq����;Hf]�	2 D��n~n2K����+.Pg�XЉ����T !d;
\��7��[:耾���
�G���R�9b�Z��smz����|6/����Ka���R���Y �� XX8�J��� ��ꅈy�u���}���	%�6�
�x`�Ӱ���E-Û�Z�{����;(I|��yU�N��5���i.��h�r�|9p+�'v���ֵ]L%Ԟ��3�įh41c�h TIii�PO����h�$����7ϳI��WAꕺ0�&C���>R��F��R,�9U�:i�^߿�M���g?E絿���w��#��E4yoģD!\7]�T7�-�<�(�1�=0���ȍ-(.���'�4֣ffa����������>0G�'K<`�(G-P�(���E}"Y�������V\*������.e�r��T�y�H�Ql�Ic	��V��i�(WF޻���=��Z�����[�y��H���D<iY�$kѾl�c�j�ȯ@E��?����^s��W��_�R�>�Y�eW(�J���%���d�QO;���������Oi�s�Ο��ӱ���L}dS�a��WHGd)F���+��䑂R��ʫ�FD�� �*��K;��@�8��la���hl��KUB���O%P��V��͸)x!ǻ/��4�r�"�pƦ��V��g� ��sɹ��ȕiA�W���;����R���w�.��ޢ%��Vi�.� �b3<S��')�����=^w|?�Cb�(�x��qL���4��4YZ�A-vv� ���)d}K0"
��t��i+�ۃ'�gsgQ���=��4]��+m*De�AU�T�7��e�.��р\��ٹu�h���G�F27���]��g��O|k�v��a~�[`�۳7A'�����k̀���-o1��21hǔ��x2/�t:C	�iR�G� 4����hL��p�M%���Ӏ��� �2.fq��ݶf��E�Dq]V�Q���q���dhE��Wl�hW��u9T�"#f�/�$ͨC�I�˴�(�n\�ع�Np:�2��fͱ��k��b��6��D����gb�h4���L�{om����2���|~}�q�yn%��rJ���

�_q�U<�s�rh��ܙ�������]�����w�"2�2O�"�o$��(J���"w�8rQ�����^��<=� ��o��r�P�҉FF���\1T"�-/���Y\r$[�v�U��+�-��oi���͗��+�,n�}Ob����h��k�Rpe�8-=݀Z�q�"ДJpX��zKҖ�Lk�

	aK�
�]�����M��E���?�+!|��Q�������z:�>\C	a��|����F�1\�[� �ߌ��\q�F�f���`�����M�	B���ke�n���j�����QJ�ѩ������Q'��zd���C`��c_+M��k�O�]����9��l�'�h�����|�s�q�k,�RO}I5gW1�QP���ƥ��Ƥ�T,(�0K�"!ʗY���uu"{���dn�d.�/|@t,\��.���
��w�gv���"�:"am˯��Q�u얯��Ă��7-y�Ѯ��4�|:��k׊�^9T��M[��9�9�h��]���<����k�VE�.��V_k�w=���s��"m��C�i�i_�o��2S�IS����י���Ɵԡ�_��V�H��5��ٰ%��n�ꥯ�Z3Y��ьށ����\��(Ϸ����f*��[���n�3'hY�����QVsD�);�M��f�<����t�2i}�4�Gr��#+f*�gT�Qc&��*?

��Xrl�%Mg����ʽ�c�,�t.4����5���� k���M�]����ў-��+;�k���g����:�}���4$7�[)��P���:��{�T�`2T{a��O�1T�x�4N��fY̩��֦��ϼ��^%�E���������<k�cF0_��A2�C89�ɉ�y���-l�ظN��1.�olnv���k��U�&�Fh�Z��`R!g���Y���`��l뼷�Γ�Ƭ6<:u��b���sJ;��=6�p%�_L۴��=�Wzyv���0:���H#bܑ���&Vֹ��4d�>E�?c�/(��DB�x/��ʽ%7|1M��&O-�U8�ƲV�A��'���&��7���ivx�Ѕ�{ 3��[�Oen���1I��'K����HK+��QUn]�]�,$���?��7E�y`���7�,����J��~�t����������͍��ŗ2��1���y����u�FC1�:�{����'��c���~5�?l*�9��!�DpL�W/)�|�N����`��Gw-Q�f�T�o$�w��ѐ
�ӧ+-���Hs�!����0���E���󎮏#�feeᇉ�`����NN�-g�]�VW?����u	�������j��0s�Cn���V�	zY�,�ޒ������3t�#�_������,݄f}������~�s������c��/:Z���y�r(��������:{����T��|��k�!&f�Ċ������m��V�~�-���.��)�U�=>u�DՋ;w� �T�F�� ��
�sL��$�흛����������oު�;�󥵛��ieF)D�8ў�'B�`��T�8/����XzP	��8����6��h�2�58u��2�
=������ݼ�u��^N���i=��w���� !�#TN�k��:ȆD��,�����MT�"T�k݄p�Uf;�X��Py�YȐE�)���(���<M��R����'-�`2 0���`��J^2Z�N֒����鹭`��W���o���X-��
!%�!**b}j�f�J36O�ut���Y��T���7p���Z��\�7���;uu�<�ǘ�>�}�"��d4$�y����[H�Q���P��ezkh��h�1��u�\��M�e��2+�Q'`�rL%7��[l��'Y�=���wp� �n̞h^����G�u�Eut��F1*c�H1�(E�� �(J�"�� RX�^ņR54�Ra�.E�^E`i"�KY`)��ܻ��|���{����w�̝)�cd��W3=�f \����JR@��F��Vr{ �ˏޞȃ�F|�_m���qZ�V�SQ�:�`L6�37ڂ���w�%u��뭇���Y��.'�bHv�-at����U��nw�W|���nrQ6)!b����ݽ�y�J"�5��&;8}����Q��P��4��Z��1Gu��9< �9� �W�c���!�D�b,A�} �b����4���].-e��-LO��0�vZ#� �o#))��2�z>�]�\K
���r� /��Wc��m7�+q�"�wpvfL�y�U؏"x�zl3ei�ee���;F[�U�U�����|��i���R{�������NAy�#OMo�����5�R,N�xX��$�^�֫>kщ���Q�Ϋ4����@T>� �Vr	�{2匈j|I R��4�r@�EH�5p;�_��
($17�nw���9�-�Dj{�~c�_��ɖM0P�ج�f��)���nt�R��y:��]s@(dW�>ή��w�}i���.*��'�F\T�j/�z�Nl�,���ܐ�+� ��	I�{�\2
��&g���0u}lsn��T�e���js���>׶?�M��[�D��8p�;�����z͸o������&��� �* [�u��7�5���9-퍁�%�SQ�DH��'��)==�x&N���:18�ޓ���ڶ�ኇ�G(����ӊ�w���������U�M~<6�ڍcQo:' �n���a�0F�6�\�;^N)7i���a�M��!�:�5����/	L:4���~���X�<�_{�-h�;�h�z�`�l��ԥ�ը�����%,�W�?��Q�cSdH�}z ��=@A�[��ňX[����S�p&"Q7+�
p�����I��Q�Z�D���xZi_�z~��%��� w<(^^�i��Fx��J  8"�f $��,��'S�ǪD���j��d`���֯�	��b�Q���0�P��?� �J�H&�E�쎂��j�_&�Ey�F���"m�ѡ=/���2�y��\.�I�#60��̏c�G2���.yt����E,�� ��(d�j
8��#�p�D16���G����`����ޱ��GL�v�W���DTk�9����?Ⱥ����1P�S/����Ťo��2�5�Y?t��x��~�mX:/�U�=x�69Jb�\�$N%�
Ċ�(B�c�4S���C���G�����l���v*Tq��T	x�*V��{�J�	�0���L�f �=T��,__|� ����,���q#v��ΐ˟^¾�on�; =
��<^Ŷ��Ch�@M:<+��*䊠��[Qa�����%�*�'�;`܌�B�ؐ��6���]t��ki�;H�9�9���z,��a�@����^���z��~z�	_P^�t^d�F t!߸����3~t ��rS���['g�V>��hv*D��BPO})t�J�m��s�P%r�(�x� -�� ��N(ŏ��q��}2+�v��%B�BK�����@X��|��?��_�K��p�%(��=�
�D/3U�h(؀�Pmv�3 :��F.@��G�s�-t�ŵ��ʵ�/0�����y� .xTe'�},e"aw�	�������������6������.��vV���!�4�L[�L�a�!��&O�nG/6�<0:���g���f�}�<��z9yoZ�2nk��F�+a|w8~G6�c6)�G�u�<�"˲�0�QQP3W\�k\N��+l��9�r�؛JK�GOgI6�F$�!�E�(���w�ϖ�2��>�� ¾�R�7��!Z���xb���*��J���HN�C�m��=4�����E>���NA>�y�MXo������ �BP7^�>~����'pѝ�6�����]]	�:k�kH�P�J�zO`�=��q�zry�����6��!��S��Z��GN�����m���D�ku�L{S�$��S�v�`8g;�1��A�7�zR�Q퓟;�����O���Kn8!�d3��E��^���s*o��������`Q�`@��G���C������#W|
85��OZ��P|4�
�c���rP��S[ےl��h=M����z.�q[� RֺT��m�o;o��F�ah0_���A��oT�:w�X[F��3o��AD��7Xz%�7
��6$�=5�R�^d ׎E���9���+q~tC��$Du�E0��
��Զ�����Ц8ަ��oTP��|�M@�D�^��CN�����5��M�w]� 2�`�g��x��ax����(�)�$�����_� �م������{�aVݾ���&�9x�"P�	��S:��VOp8�̃����WIT��C�˲yqd�Q����\^7e�H�E��[ͬ@���ӥ���wN�3�;A�c6���mb*�۔TO�@ �������}^�fSU�LDe�cy����={G,�� ��c����I� �[r�1�n��9Iϰx����*�8�]��.�q]�	�|xR�c\��A�3��׬���2���V�N>�F?#���c�06��!��j�����c�ZA��{�G��!ѐ/Ҡc$���U��m,4
�����=�¿�h��34!�"��'��P�P���e���#������������q�$�W�2�.^�:��	ňXR������f���^�[*#�����	S�� &)2���/ρxF1��F�� ~�M7�Gg��n��x�mj���&"�sbGs�}����*���߶M�%,z7��5�)�W1�X�>]d�3�.���Q=%?�J�; ��p�"�[�\|Z�p��#�F�l'�+����xӥD�r�@��S!��A���]��czR��DJoQ���َGٸ=[����|ja�-�C��D��� ���W"�3�2:�5��c��3$ :=á�j�� �3��Մ�g��@���b(�LԶ�<=����ٸ�%�Bȓ��[�tZ��&�*���DoonN�}��b��!)���c�� �6���0|�����V,�O[G���X�}�Y�S�b��	���{7�6�Ю�8�cF����»�l,ԍ���t?`v�����G�'�A���Ui���e,��`*\E��<�@��/�;>j�PN,�4~H�SV����dC>}�]B �M��R�Wru�	x\�Z�Z�F�@��c%�E�UP~��F�a��:�����Uos� �P-? C��S~�C��l\�(�h�y�ײC |Oڱ���mA�n���x�>&����%�y@�Y��}	��A=݌����a��9n�����'�'�6�i�&2�����V����47�l���a5�̈́��D�;��#�����y�I]6Ρ��$�����F����x!��w���S���0�4������)�/�qd�N�FJ_� ހ���s�m���XL{� cZ�qy�+�/�"�VJ��}s����MT/���	��v�4
1�q5��t�8��vOJ��~��Y$*&5��A8��I����P�������)}��j|�[��ST�ȿ� ��D�@[hQ�� �c
(~Xh��&? �M�?�$C�!����&ئ-�혗(���V�r�j]��\๼��Z����Y�,�B�6�!T�Wb�~�8Gao�n2Aױ�ǧ$��ۭ����Ș�/���n�-cv8�s�h��J�����������Rj�l��C��/*���>�;ji�j�>����I��M (*n�+/��GV�����^���.��5v������^f_��A`x�G�%[��v��=�Ї�1|[bX10�.�ur�Z
rJ` �ʫX��K��������i�8�rA�: C'��D���*RT2�#��kk;�\��ޜ\-������U1�'8m�����ѨY3���}rH&�N@&Ƹd����`NW*>P�'��$
e�urU��mRz�t��:u��C*F��a<���s��m�:��#z	�^b :#���dol��h	����:8����~�J����a0��V9]�+��2y�4#�Ţ,��Y�$��[A���	�Z�����4a���kA�������B���33ڮ��/��"�h+Ȭ4��w��W��x�mwP�v�|�'��a��f����BxU��p+��NN	�d����Fp{X��)�����q4�bbx��~(�����P~,74�Ȓ�"�q-�r(�z�r�OS9��h]J����g�iOY}�O��Xբ��U'��ɳ����2�0����F�<%��1�����Y۬y	�#&s-�ຓ0Ћ��}6��t��9�1�������C�W�6n�"y냱Z�qۤg#H�  Ɯ����Yn���`�2+��� S��3�bj.��d�B���f�z��7al��>=���b��(��Pu��"M�o�	�μa��RTq��*o�vOG��妍���"��NM,�?��ۯ�EׯJ�6@����
`3a�`{#���ް�l�| ��ڳޛ�u!*�ʣ'�h�p��1ٲ��A8��]X9v�4.놧�j@�Y�΅�Fο���Wu����]	�6���X���VS�T(��ܧ�����Y�N���m�C�~L�߂�%�%Zo��H����H��L�dX�ķ8K���}7�n�C���\�k^�]�y�mр�>|�X��(&+�H�� �P~���|k6�׋����
�>�ᬄ�م.����>[�:]0�4n.d��k���F=���%�����	�X0�!N��8|-*��nY"�Lfe�/T��٦�!թ	�'�&g~!���}�J��8ݎg!�o� =���`J6涖�.�1�C��eC/�(gi�|�Ri����z�ꉻ��o����d�+|���o�	"6�L��(�̻����J[���^\��"��wo"�
O�R���˧x���``�i�bY�Џ��r�^x{��
H��[ȃH����	xC�k�e��v-�r@2��t�|�M�~�����i���q��on��t�oY�,��~�睅�8���H���L ��?Ru�@Ner����6��2V��#�&t�� ��j�B�O�С��"�)2�˧�5�e�B�ʳ(l��ͯdc���,�����;v���o�,��k/��6y��B��0}���~`9%��In?h"fU�@f&:�2���L�4�z�������h��&�%<�����\����*�!`T�Ȩ��	YD��#xL�B��yc��gv焴"��+h��zr�V���`����
�[u.���l��+�
?w�̷�̫Vb�
Jq
��MK����ծI������F�O�iH (�MH`���r3L�:wS:S~f �jC7^����A� {��q��PJ�f�����|ł���;�a��w�c��a�� ��J��R��[	��W�(�F���6��.{.��F����n>Xh�M˥�)�C�1�f�� rVrr �[B�AM[\XN���R� 1	��i�oy}7���Y��Nt;Gx�I�õ��m�����g�>�lh���� 6TI���ۍ�Ehu�7D0�����;��"v*����B"��)�5������	&��+,���{9q/I3�����އ�/��V`��6a��@r5_O˭��I}�{�n�^�@�_�<�Zxj�R��N�������(���}�]�<6Qu}�~�����c�D=�Ѐ�8{]�l،�/"���X��z�P2����h	Ovv0	�q;L�ݥ;W�F)9s������]?�{���&��^+�2.'+����¢ʁ��-oz�})Q�WJ����׬��/�F��2e�4&V�FO�f��'M7%\0�d��ؔ�ed�6�誂�cOS�a<���]9�XJ�T�x^*/ ��d/�
����t�b��ls���6�g6i�;��"�y'��Յ�=^�$�fp����v����ۧ�`�L)��hbd@���ꮔ�E�5�e�j/q.�V��Pd@���a��8�mr%UTWl��$�D��������F�]X�x
�R&$��z�X�����$Dૼ@ �~6x(߹���c�(���f5ɻQVm��!�(T���"zc]o,��������&R��b�zϲ�U��D��Y��Z��К~�ng�FS�S�����+���(���&��F��8�%:��q�K�.ho�V�������\	�O:�����6�x��Z"�+((�KӀ�J��h��Ou��>�<r�"j��=khcʣK��S.(�FG��������+��n�۰�8��zԵ	�]�y�����Znn��j��-�[.�jw�F�eN}(������WυwD;,��g͉�+s��5�H[�#���WB����!1�{��/#:�L�9��c���i���fz���n%s��o$�������m��=��.%腣n�S���-�ߕ���>���@/l��]�j�<l����;x?%V���$m�z��]m�)խ6yPtD�S{���{��&�9�1M����t�G`�,Y�1%��؋/S�Y(jJx��[|.I��_c*��w#C�� ��b\jʶm�[��`I�N�������N3�����h��Ѱ>�);9}�2xכ�[�n��L���T��������m�pJ�Q��4>t�����iW�u���Zp����e�O�>o	��;����>�*�I�'c��tf�{�>��H�����n�|��w��������/^����^Y�.�	[+q���41uV���(c6ЯVJ>�u�\��8\6m�Y}#���۲�F��%�֭�����"��5�[5� 81.~0��t*]}��낞K�J�dk���$*�8�;<{8H��KDҗ&�i�N�n�q��Q;n����q���gQ�aF>����i��$�<��ކ��l�./��N�;]��~e�:��Ʊy�����𳌇	^�y�_��4�I5V���u����8�=�T�mQ�U=gN=CY�\F��&H+&Z�%[��YSq�zd���/t�����ꗹ�0�O�����k�~�.�;oE�٣,`�p�C����}ʞ�!��4/Mt�4!�[j�&j����CC�?G�
~���Qd�e�z�))�<",.���C�1�-@=���#�����Y��*�"�H�c ��ܶm(ى��0@��"�T؅6�0¬����:$�y��q��>��,ا-q��ˮH��f����z8qdC;]ch����!i�Q��@�qg�YCBB���f�̧�A��#�s��u{��@8m��z�#�&(p7�|�t�]����� K���=��H+hÌ�!M��2,�x����g����I���2ܶw�OP??���>��U'�c��f��Ð ~b^��Ky6
?�P�y���)�{�,�UkƤ� e� ��5��.�|��+zj�MY�hw��|������,�z��Q�!����s4������W��.(�]���KS�˟�7�v_�f��o2�f�T����%ϻ�Axo-�$��.Ι�n�-s�"�/M�e;L��ͦ���+A��L�ժBDAT{U���`
RK�:�����P{^E���7ڥ��(}Y>`դ��^�'W����Z�e�`��r�������ǵ��A��6�&��`������H��!J檞S�z�&vL��^9�&w��J��؛���)�FOO�,����ƥ%+�eJ�����g��Oc�q��;|C���|�2N��o,e-��3<�܆�����#���:�����r��J����B����T0���O�u|�
a�\�|vM]����x��˶�]1�'V�%(��Y*A��ʕ���n�%b���v�^}�9�ZY�Z�����?�#;�W2�G�@#5`�`�4'�/[a�O�Թs�w�Ǐq��W�h��#���$7��7�j��	�} 5���VO6��N9�`�m���N���32����vl���˗|Td.;w�����^��<읱�r��:���OXT-V���--߾]u�}�8�}?E���
�y痧��~��-�?,�D��C�`�=x35R-� ɇ�ŚJ�Bl1/%녇��x��ִ�����U�/����o�y���"'��^8���?�����f4��<7�~8v�3L8��r��.S�~[QJi�{��K�ю~θ���s��0��~�0h��B*J�*2�p������.Qڇ�o�a��z�:!**2�o�����Ń�ū�2/���.�߂?�=�2U�2qc����n����DU��-��ƤܥpR��*�n^1A����Oo�j9���W�^{m�n`iްM������s
K����G7��*�4ͽ9���K" Tg�|	ʑ�6YY�˱�[�;���h���Q�9�k<@����d�u��҄5n%���ƻ(��mch���h�p`�9�����Q9�LA[q�e(���O�epO2A��0!n�f��8~p����[��P� � �A��)(�>��o������=N2��"�/���Ԥ�ƅu��M�́O%Gy�ρ�5__��<Vd�溷��>\ER׷)�J3ٝ�Ln�m� /+�/N��#��A�qV�R�%$߇]$GJ�7Cl���<���h��<��B��
��{��u½|�g�j������u�w��X�1��_�F!x}��[�z�����K̞�: �y�" �A��ƚ��@v�JV�w��+',� Y �yfD�!@@����-/���l�
v�F��<���VnJ�r�({��B���C3���Q��o#A���J���������X��엡ܦ̓�䚹9�Pu��i��˗A�tt�ݗ��C��1�:J=[���ш��Q"���:���N��E�$��6�j�xe�����2��Q��>J��	��/���7͇�q����@i����O"+����oHQA�#�����7��/��U.1(YJp(V�l��]��G��!b���3Z��W�a�:��	�C��.
����_��������guu5$�P�֥����qL0f7��8ߵZ)(���O�̳���P+���vx��ƕm�x�L%M����fR��&��D�xȡ\y>���KzO). �Y�z���N�z��ϟ@Q+3�A�B��\t4�V��n�r��'f#���]~B�~DP�A�8����!�K;E. �h�u��&�Ck�����[%7�j�ع?c�Ƙ���zf�3�x>A�g�V-Ŕ s �o���\/�)�p����?��Ck�z���=��̒���ȓ=��OIC���f\�7?ko׋-�U̏e�|o��U�tm欤, dv��;�D��c:hL����	L�;�B֓�C��1�L���%m~�ing'ũv�!�˿���@v|�e���Ok�u!��9z��xez��h�JxD0�Mz�.�u�wƱ�ޡ¼۴V�,���p{N3�􃠒ݻ\{{8{�r�Նz��eo��8�;��e�Z����[�2o_���Lq�\m���"��U-4�I�ݞ`j�S�8����m�����is�֜��g=n����S���7y����m�G�2��&���ՙ"�K��)���?�n@�W���ya�7��B+ֻ�KWG'{��� .���DA_���[����O4�< $���2O��#���-Ŵ���J�k#zR\S�r������O�78�Q�)��	� i6�(�2�`J<���Vn\���=2�8��7Q�#cc�a��"1����{Z��,�Î%�H-��T�j�#������|VN�s�����=�w��ۅ��֌�LԽB_8��NvL��<��+��;�!�;'��]Lj��}�,� ���a��R�R0Hy�}��maX+7�r�[h+�,rw���Q��{��nY�.0ԁ��|LNQ+�N�c�׬�.��i{{;�EPq�A���W��CqO��������{t�8��˱��kv!��P�hZ{�g0�kB�*�&oNu�y��� _�.�Ր7���SX�����Լd���_��r�HuR+돷d��	>�2�ڡ����57Q��$�<F�@&7o!4C&SM�Ug�����f�.�Ⳍ�P�ڊF����7��CFq���9���e���9qD}Kx{i���[�{�\�C��"����~W$�Kʷ򅷓!���\���*6['#��}���;lZ�ӨSJP��N����X�y^�&+�QɈ�f��@�^\�"*�7�q<����wl�B^����Ug\�: {�ŀ�{(8�L-bv�:�"*'�����LE=����2'Yށ<U*�:8سs&�	���/��S�0u��鑎�N�4��;��+˯�q<8���R�T�mڀ����R��e�J�C�>5�D/��;���:e����hy��0{�:գ��Pٻ���]� ���p��5wsC���]cR`'��`_�l�����;����;�ĝ������L:Ȇ��G{e��j�_���9�d�^TP4�<��r�I��aC.:���u�6�l�g�W�K*t�RT���v#M��1c�h)�<�p�d��k����0��R����'�,&�!Vc��F��a�\��&�Sa4Lk�]6⎅]��|�47I��:��i��UPל�y�w����];d���4��L�8���Cc����D�Au�ڧv��/R�&�X�J붞�l�L�t�P����%XB�l���(������+)�uJ��D5�bf���SB��K7�ߺ�n�7������ݿ;�Y裭�JroW�Ā�Aŉ�&������KWg�ȆU7��'�*n!��:<ِ��yG�㬴��N����7���S8r"g��*��M-LtB����WPJb���OZ[�����Fљ �ߵ ���|���w�R�}<�~t�
�8C���4�=q�h�pP-5u6 ���[��ؼ�E�[�PPV'�bH0�Q��R�=mȱ���3P��D1-p��� �ݟ�r�WW�����%K�v+�X�z�:10�6<� ����$J�*��8�ʆc&�ݔ�#��1hX
���"�Tr0�y�a�6��f��r&a��� f|��`c��VE�X!�۴n9�95eo��_����$� HCb�?�sB��Q�.N<��;%�dw���d9���o�1�nNY-�i�w轢�o�A�OE��=����F��k]�r��<����� ��N��q�.=�u��l��YB�ؗuho;�~eks�*�F�J��2q4 U�5'G�&���N���b%�3{Z�~�r������4~DE�-yX��������- {dd��hz{�D!0�w�l��L�q���~'_�_YA�Ǿy����'�U��Ӛ�/:&6�vȏX礆�'�.�'KWMPL�g� ��'�J�F���e}����㊡�څ~������3 ���x�n��Zr��Lo��OY�@��Xz̷6��4�$�] �&��
@��+��&��Ç��e�l����7��gfϞp+��Rl�dl.��R�I�wZ|��������31(�ʋ�;���5�"_�D.i��w���#
� ����f�����]�I��_P��:��xnC�o��?�Ր��rAy�"�W���ݧw���W��|��!" ��%"֕*�m��L���W�7b� �)��ĺ����.���- a�蜑j��n�zDn&_,E�3_��l�v�tu�Z�,*|��s���@�5k�C5�]/A��(�U:~QT5��9�)����㰌|Z�60Z�%JȠqWN|��T@�? Z�;�8{��K�577����UjQK��U���/J����t@I�UN��V�%qz���)�� ��(8Y���F��..y���<� �ğWe�׃<.�(�M�%' Dv+$�p&j�����r�5�MZ|"�(:dȝ~�e�/rl#��H	�����0�+�f���&���.��CՊ�5�Vko�Cc�+3�Hy)�{��P}]��h�R�b�j��.���/\#��I�>��j�bd������#��@^',K������㦓qg�l���_�Fڃ�O�F� �����luT��O4X(�es���b�Rz�K꺛;lӨ�E�"���|ʸ��(�#V|����[=v���Z�-��۴Jx����E~K���e8�\�{;�g]��c���Xeݠ:i��_�	7Y���D��:�H"�d5${v����[=��xų�m�kЛ��s�m�1_dL�*����f9 ���\�(ˍ<J~f��띜W�ٿ�*�oF���oP����4ǧbګ�����鍊WL�ԸB%��p3�_x8�����q����x�fF��{�8���ݘL�=�Zy6�VRd\��!2�i߫�\7V�ekM�|ƣ!�2�b�^��T��[�tUu�� �TF3��<��{۽�r�]W�?)=Ǿ�wdⳡC��W�k�p��ʃY��e:$�6���[]1��?P�������i��.��X:�} �
�^}tN�O�7��O>fg�'���؂52���4+�b�!S�x��z�/� m�=Կ�d�)�;�' ������$��^�q=�^?�!A֞ȒL�l�ך�ܷv�%ߜ�;�x�/UM��e���̃x(��(w�)�' �6��� M��&��Qm��Ǘ�[��U��Y��Lʞ����'**���v��k`n Z$����T�ou�G������>��g���#ܭ:)r�V)�vS�G���Hާ��)���+�,S3ԫ9�m���^�쾱� �<��wCnl�͏�K:�����BO��y�#r���@ x�G4cҿ��KoU�M�(���@�x����`rt}�ۭٹ��L���c�0��N��R��k�P2�\@$>�hv�4w]�B$�������!��ׄ���&��m &�6Qsj�0N8���<�89M�'L�i�g��1/<x8L��B�/�� �QP�:T��@֫!�q����W�Ѧ��n���5nP��շ�T�e�K���� P��-��3|d�/n�1C�<b���p5B�ox�?��.#�:�7'�O[P�{�K�!�F�s����d�0X�4�4n�F�����S�Es��d�Yy� m A�����m #��x2죈:��YkE�l��Y򶟣r�c4�N�j�ơ�0܍(U�b�@�:be=�8 km7~��a����z?ȧp���	L�qBF����k�(� G�fK-��Afhj_�'Yq�LoP �=c� 2����&KS��2�*�{��������M�	0��T��0��Ғ�� �\�46�פ�a�8���|R�a��mb��2Rjr6S
��o�)�_��Ю�TtH�������-�mp=�ybH�\ ��7�+UAa�`@���n���	�i�w�F�Ͱ�O8�����[��h葻���E�^_$�����ט��^: �rJ�Y�SG����rN|��R�C����w� �j3[4i�IU��ܞB�GDh��E["��V�|�_Je�A�Xt�%�͚u���9
�|_��`�Q��&j���-�NfI����'����^��$��@��w=�K֍��S��_�,��3�6���u|��a{�'�}�u��ѻ�e�̉<b�1C(b��s�m6>2[�Vil�_M��9��	<\*Cy��gUP�d��@�Z��^|yni:��j7'�i`��|R̷ɋ�\�@	$��Ʀ���X�o�K
�Lej����OS��1��y�X�E#,>��y���Zh��O[[[�|t�ʖ�zĩ�o�;��7���ʔ��zES�?j���#���z��}��\F�]��L��FY*/�G����� ڂj�$==���SP:G�G�������ny��7R�K����M��W��V� ����N����C:yS�<wG$_�Z)Tn������"������Mn5Q̗F���wl�"5�����(�^kd�����70B��qZ�ܲ�a�T4�)���2:��rj$�KB��>��/
ܡ��4u��F՛����/o���go�O�9 �T>��A����i��U�8Sp��0��iW�;��_��y��~8|�A5�l��8	��'�)���s��Nj�ڍ���|�SF�s�Mޥ��'���<n0[��N­����!�uZ����1���(�e��c��+�(|R����J[�������yൈ�J/�8;��ZZ���m��p�68hG��3u��@��0�	�E2$[�I&�׉�g�q�4(3j;���Y@ПVW��=�
�h`&�B��
����D��l?�]X���G��{��
��T�*Z�=�d����WN����e�t������rQ�|~r"1�Loy4��Dz�4�Ɵ�{��_I~T9�/:�疝0+Ss��`g�Ǐ�q�݂�a�@�U�@��?�JCí�x���1��r\Z�za�Z(��E�����L����%�̠�Fض-9Cv��փ�_)�oLZY6t�2\yd��1T��F���XH$�.��k}�c����[ԮK}<���ԤYuS�;��-�9�
�#��m��j�;p�۴�R�&q!m�Q���<
S[��*N�ӊAx�Li~�-�*�{��O^��~�\�Fa��O�&��� �a� ;t�CU7��5w��91{t�fB\B�K۔5/��1)p�����w{�6�����Jg`��^iud���Fݶ��R��3}hJ�%AOl@�介�S�ܜ�����Ef��7�L����J�B�P.e��Õ^ �;P���B�CIm���se��Z72��!������"�'Y�6�[`��rs}m��V�n`/���"v���]�U��Y��xm��(�h\4}::S�>j����9�Id��(���i(Ń`:00 ��
�W�/�_����'��{S���y�Ά��{̔�����qބ�����`�r��>D�q���e%29h��^�a�:�q3j����ԯ�V�xv����+�����P��e~(���:�b��˦ nɆn���������b��뺷�ˤ�$�j}}s��DS�
�+�f�}��q��p���c#��\r^��viD����S�����&��A��T4;�Cm���A}�x�����߰딨�F6Lb1_���y�}DͶ-�GK�¶I K���v�"0�@�G�PBSE���T.�	n��.mRt-$G �j䩟U�ޑs��������7�9ܭx�<Z��m��A�^Sw�_,s��'�-��F�i��@e�m[�Fx䱟�L�g�s��s�<���r� ���B�q?���w���M�6��#��/h����� �`G�N��=54y��������M��Aզ���g|�z�c����%Wd�I��3�h` P=ؔ!n����_��)TZ���P@���v���,Lt\�<.��w�����f�
+׹aq�|���z����[:b�3��R����F�9��)���Q��őZ�A�;� �(,8g�~Ě�CKV�I�yN�p�����^Ya�Ǩ}Fjx{{��f%j�����H��z���A2��&pK��D�+í̋��]���¦&r�k�P9hR" �j�T"W�����֞%鑐�?Ev�.e��s�5�ޅ�ل��-7
c5U0�6�m�ݺvݚU���{u���������9SC�g�	��r�(X������Xxb�t�;A��+�b%�f.���N��q�g��T��<�*��&**)e�<��+P<'��x4�f�N)�������3���@�I=}���m�f�۟_�ȟ��CG�����7�d�uW���-����",�S��G���9��/i l<�GTDD��62���y}�wѶl�!�.kKC��7����
��_���N�Ww[��+z��q��#���'�J���� �Qj)���C�޲RW,B�׎G������^\~�*>Y�*�zo>��u
��-������K�0dＯ��+��W��M7��.�_D?+��z#^FG@�r��r�����9z��nSS�v�S�bRW����g!Pb��L+�).u�6��K�=x�D�7��4n��P�k��=E�����jF�#�ժ��$�=��ސ��#�d��oViT%�]`�xC�RzkU�Ű�l�M�tN)QF"��٢�?�b��e��놮����?�rA�/0���hd�?}d�A ����s�U�$h߆$s�im���sB�c�⩆�S��J<����AHs��kR�㭳���֖'��Go�u�ͻ�C7�|7�<��u��FQQ1AG���	���KU�(8fl������B��*U�![���)[D�����~�f���E�MU�����l/��L�^�G��y��%t�]<����)_���,��0�޵�F�;�Qq�En��::YP\�mc�<y033�lRg�I��Of�`�pO��³_�X��@�����M)�8PI��U��NB��9��Ř8%C��v�yaX�6�f`@���Sn�/��NjpO8�X���X����}a]�=/ܐ����m�����ݫF�ۼR".y|�����o�2(
�Ğ������@�ߛ�1;��^#�D)���%[�EV�漩�K@?�G�vk�dK����{�5�;?��j#�a}�Ő������C1�t)#rssӥd~HI����.��y�:�>�_g���%f���.�v������~#��A�~�-#��pC���x�\�2��� ��yK,�<��*0�W��B�D�w��K*�;�ϻG�>�r-���<	�AQ˙[֯:o��;Ք��W�1��5wAc�5 ���k��kwq��rny&)�4�#�xS�0�)��k"�;�nu�$�
���e�����ζ����g�l�4
\ťL{�M��9������E�/�*���b�cR����[1v�Z����*�|�w�ؘ���>K�����u}_&�*��w�jxxx�ٮ;�/?ž?(ix�n�`w~H��_�����Jd��C7>h|�Q�jr�4G�Aː������Ðf< �|��x�����q�#$�<���b-�@��U{���&�g��'�Q����X������D��;'���4��K
F���R[M��hgx�s��u1�F��,��7�X/z�]�
d˧jP4
Xg�.��𐮨�D��"oι��V/={�Iq lޏ��:���&���/�0}�_ж��� �e�+��-��6\����X$:�s�-z��#����&��L���hV��fo���>R�h�%��Ee[�0�����D��*L�۹�q��:gay\Ո��n&3��S1d��b|彾6~�J`,x�ȅ}]6_v����ʴ������5u_�
.6@ GWI�A*Z���9@Y`�Df���s��1��ͯ���v*l�#�໘H��]jU�;B�V�Ɓ��UMyo�,r��Ï����@6nb��㮱k�Nj
�S�S!>&nY�����{_Pt)�mS�3��o-.��7-�E��k��q�Prr2������u@��$�Ҍ+_��M/���@6��\鳐̇���z�އ�W>�`�Z��7�?�4���YΦ�Z÷�.]�"]3�5�����]�6�6x ��PUx U�W֝�O�<�X��2��f���2.oXS��Q)O~ ���FKk�gec�D���v��9����C�1�c�`�{�ۦ/�D|��+��*kf�B�(� ؒx�<��̘�:��*�W�#?R2	�tx��zɯ�˄�=oo��Ĩ�����4tIv���1ј�C,��X��~{�\�s����1�@���v�����ݟ`^t4Ee��G~�n���ZU��۪f����rt�3)�q�e3@w0@ � �ן����FE]�T6��͜��� �]aQY�Rr��I��7RŻ]x�k�eA�q�<F�zP���!A҇��t�;�t��r�����:�i���l�u?�!��b����ɋ��� r��ҏ�=�0ԗ�O�WuR�^&zE/87��>,�&+��c>~W>"�5@X����=,��~�ر��W�~	620!�.@�M7�O�X�胸ۊ���E�^�WOpe��<	>'>u�<T5�5me�'%�K:<��2�����H�&dÕ�<�/Ͻwp:ɧ���~�B� t�BQ�U)��~�RO������1!##�����x�m���&�$�yP�ytE��W�#�}$��~�Э}O` b�B��h�5�ҩ�`����*����G����O���o�T�AH�DM��¯�� GӅ�;��i�����_��4�L�@��?����{���0�����H陪LJ������m^$m����(�(�������Ϡ�_	
v��ߏ�||4�2�i7�#�*�T���#eZ�ݗBg[4+��~E�u���?�;M��`��m5v�Qɟc�6`u��m�ԉNt���:į��t��]e+z�)t�i� *�1�3 �s1s�j��09�&�B����0XP@Q)��=��N��%u���w�g� 	j���w�n'�;�X%�ߎU#��������K���f��mn��t��ټs��v��J%�I� �y�$\���[�uc�b,��5[��4�2���t�/���~�Qq�f�y��ɖsF20BFa�'j�
J���iMew�%��6�w�զ�\K�1=��/[�Z�K9d=$�Sq�k� �bc��. �D��.�l�މ콹���˻ޭ	R�5�������{�3�:LR8yO%R�Vz��r����g	�	�#Wa�rk�^�ZH�W;Rs�`�~b�`n��	�[۵�
2��uF;�X��V��;���E�Ʊ�nǑ��|7����Kn4�0qx�2�
3�һl*H��8p"��#T�L��\[G�Є2��^�3Sz�hhz4}�s��8�!��!��=ExNЪi�dG�K�r=����1 7Nv����H@��uu��� ڍT�!&���ݏ/�za�T�q����u�&���9���x��CR���r ��ҥn��][С�|0��b�&�n�Owv��Kъ<i�
��C�lV4�_��nY��u�p~�10��v�L�P�Щ���q��n!�?D�@8��1�R�N���Ӱ�����P�@޷�����M9��]T2t���]Q�o��'z��,e��$x�6"���ͼ����K�{R���^��c 5�6��W����A�������M]�j�[�-7�W7N��F�j�Dj�{^�J��s��f�䬭KV��6��\v�ҥ.2D�	�Ni;>m#�L?I�9��nyOCHtPKu7)_��J_��9qFS�fF� DPċo[���v�)��9�N*�ZTWQQ����c��t�%�,��?�K*��v�%>�]-�E��{�s�L�l���w�0{۞���k��u�w)�˜�Ka�/37�8n�����_Ż  �{������^ߊG��եP��Y��Y�}nV�	��˽{�{���5��3��/�S\y1�����b�N�0E�2%���ۏ` y#��PT곑���HIA�4ȗu_�${�yy/� t�m�ked��I������jr�o:�JYY�'N�9Ȇ`�/B�>#��ư��p%|�x��Q��qYf[��p�����R*�*H�c�"!! ���� ݠ�`Q�H����t)!"% �t>R�����~���}��Z׺�����w{��ğb�/!3(�4L�J�rq@��Ò�,��YN�/��8��~P��+*��R�S���>������#���C;��ɂ+Fp��YN�b�@�U����.�]��0���f�$d��C��i||y��Z��`+ *�W �og`\u���}=_F������y3u����^����f�v��ϼ�V��Q�ٹ_=d#r��|d�BO/	��Z����$�' ��}�\���mJ\�A���&5U���9A��D���)*)]?�3ښ����tt�Ed	g �	�<
�B�ɦ釩�zƿ��6e`�Zp�á4���.�i|o���r�#]tf���uDx�F��8�\d���,L�P�Y�eA�ys�~��Ă�!^<�����է��n2n%���g��y��(��q�������k#���F!�i���a
����I~���*�U�.R>^��D?)� d��o�GK��aѹ�?+��dd���}���١i־Z�il�X��q�Nq\��'�"�j�����d�Za����I!�N���!���|����cB4VWm����Y;ͅh#�Ј+!��y��`~�Ҝ;u��C�օ�n2v��`�c �I	G��*[���c�?>]������~w�r쏍�8?�9P|��l_7�caL���.e��o1��hEj'0�$%���?N�/Q�W�A���2�
�
�:ζ��^�&(s�MʾfǬ�Q��]k�lԳ$vxK��9=SZ���Ņvj�q�#A �����db?����l�%��^U���&f%��+��x�a)��+n�cw����jq��f�9���ȱ8aINi� �:���=�������Ǐ�4�2vX��>���m�(���R����F�T��|pآ�c��<�\�3�5�<�M<��yR�M��|n���~_�����ʺ��%y@�ǫt�`e�T��k-���( GL
JB�&�ivL~�	:�k�vK�k.�^^�13�t�-e����Vd�^�.B�����4`"<�]��)���!(x��) ,5y*NB�9R���!��e͉�[L]��|��y�ӑ���滪$Wڠ�x�%��{��Hy��?-��V����u�Gz���_L����WڟO,NV�ʘ�౐J�sC�>x�ZPJ�hct9��fmm��f�� =�Ԡi�]�o-"�r��R����ț�'=�����VS��(i�H�E��[:L�����_��@�;L�c"�t2@��Б�����_�_`U�wv����ؔ��J�����<W%(h�U��]�����H̛_Y���$ux�ή�������/mY�ب��p�f������>=>HpJ�q(6��H�(�Xk7�V5f��l�P�Ԋ9`!�CBC�(i���̆��+O��f�h-��v1���]�9`ЛfW��L�#�\S�Y��]r��!��fO��d�;��|b�u�l�UEGGwg��WTq�A���hg9福���6��=_r��5<
�&>�9l����S.��g��D$�T�E.t�t����p\!���hcŢ,xO�R�b����܉@���Ts3��7Р
��V�M�#���Ę٘f��&K��^�4�k��۷��3Z�;"��즳�gk����m���ϕ��8�ɢ�4�b�����0��?��qX���uKk�9��!�Q1C\&J�`� �ņ9�ք����ރ���{� @��p�Q>�F��GHw�Y+
,������/4QSX�k?arD҈[��qa�='��G/��5����HT�O���y�\�\��p�` RJSEq"��Ȥ<j$5�|��"�{��o���wwR4�N�P(/���prFdoYr��$g�y����α��a1�`�G����j-D�)r�[���sK�T�����LWs����z��4@+��mK/���Z��k[���F��@S���H[��dd��������s�/��ݝ����,>ZX|=���̯�2O%H�CNW��*(�AHb���0�����F�Q:��2B
0%e%O��q����I�݊aFFF���+�ǣh� ��ўc�封E�����i+ݨ�ݱx¶��yp0���篸�j#�Q�Q{s�rᜆ	M/�'�.:^}�l���ʶ,�cslsBn�(�:�-�2U�L��K�ؒ2?��������8�m p�������.�꩝�����M����\�4�;6	kn99�!y�M"��S�\W��*�@@�9�o�///���{��D�`��DV��� �
��~�r,j�Z>>��m#ZePvD���,)��/����3t���0�E]$��;A)f;��K���fJRCva*�I�����|@̑����w9@l�v�{�,�^�=�88�K�en�ΰ|F���'�@�"ɲ��%�Q��7?�����Nေ�ѻ`��og|�N^bۯ~5���He��>lt��oNnk��V�m�=�\����R��@�'W�����UHт�r�|����}��]��옃K?�޿	���H���L��?�;EH5ygD�j���f`^��r�����I� ��uʯ��؏瑴r��,*e��I�l�a�6�nл�+v��46+&]��1@>q��Jڍ��v ;H.����Oԓ�6��I���~u�F��h���4o��+��il5M�f�u�"K
@4�xWS�a?&G!�X����m5�ZZ�������U���)���[x��m?׀ڍr��Ò���7У��|eh��TD��u�۩�g���L ���)�ݛ��o�iʥ,Q/'Qk�ٽ�E�CfN�N��-!YV�J��9F �t��/�$��ʲ��eJ�~xz�S5,��y��C��yh��ڰ$�dG�������0���j�\�IB�ל��tD{�k��H��UR2�Wh���-B���ùB�9��"6�;�d-s�,Yrs>�"-О��!}?��3�+�/�!H8�f>r.���w�̷��p|� ��v�X�������L�"_���B��;�v$������{�<�2ov�O[�"�����f&��{?�Dه����q��2�ha�4�ITc��N�k�]EoL�/P�A�bd�n�r�q�F��	��#�����l���/\����Of��l�)�� d��ȯ��A%�-y55��u��u�u�;��S�1V:�yO�9)��EeFd>\��Fz�,�b�x%_��<���wfH����|�h��3��0&ܑ7��H��l��`_?/ʷy�Y��Jx���2/cs����,I��9�E*�J�I�E_����� 
ncc���KI���������y`L��^��IW�L���}/by*F��4�l��g��S%����<�g���CJ3O�[Z��5��$h��:LV�Ի�W���|�tX2Һe�늡Cs����c��-yw%��,26E�:�0Ҝ�
��7��;*�	�wOyG=�!� k��OxY�-N�^ݦfP:?|���c[�QՔ�w�i������1B߂`ZmWD�C
#-=���ѯ�֓f�#�4j�Ә�~��&0�2$jd���"<�ԑ�d��I�^t�Z?�\G����q'3�e�*�uk��u��*E;=�N�6��t�����d�JnC
^��Lz�+7ė�����I��<=-e[��CǸ� �R���^ W!�V	feOpc����v̚ۂh\,��%�ڄPOz[��d�yaF�X�����	�zVSy&���ҝ#��gee6o+�-i����`_��ƽ�b���wwfC��������������o$m���X�Հ��ҥ,�Tn��')��I���Tr���&���ÝƲ��cR����hhtk�{���(����~ץ����C�ny{R=[=^=�\8�T	�����n�L]Ĳ0V��ba�Q���2�_ř˟���Ӛ�F�c$�Z�mLm??���DL����of=]E�a�U��09]��0F�Exz��n��ݘ��]�Fܳ�X��[9]�Wְ�����4��pC �YDh>�]_�XN��q3']7�`�옷�d�U���za�����con��Gޡ,p+�b%)���{�|����(5��ח�4S��G���c:?�p3��=���@��I1�y��f�j�?�8�$w7l���}+��}��G"�`M{]�E�cܛ4�
:�L3��L�P�A�q`b)�>.޷�a��Vk:S��\B�(Uܡ�E�DT���م�A����xn���Y�iۮY!���T~�>������	X�x��\͞�*��b{�!�z��!D��u�<} P����Z�;�-�*o#��#\���/k����ܘ�Z�!�X�*�GqY/aʑ'X-�x�.)'���?����Zy��,Xj-�f�L&u�ؑ	,J�F���	ׅ��c���
@4="u����p��x�ߎh���Ǉe��r7�s���ܫ��&��$a���1f����.Ї�UZ����{�ßo!��q[�u�Ѯ<���s���u��=s��
���NW-Q�݃F6�A��r�FF�6<ɪ.���߷۳�����i��VZޝ�p���M�Mm �/��Z%���?AA��}#�Wԛ���H�Y)`d�v�+��ӽ�N`/�p6h���ٔY.����u�b�r����KY�A���Ʋ�P�����.�m!�+}�$�h7��ܨ���9XៀqX}��kcN +�'���z�d��1X!��k���m�<��:PWoc��4�g���N�y����̡��9�k�$]�7���#Uv����m�j\W�^��,�JE`��Q�T�oW��A,���'�|=��'��ChRK�denњ���8� �]`a=�1��:������̗����������k߃�ۏe��a*�'���U�^��9�g?��Q�>aR�b�XYYy�[e;]f�M�w�ߑ~B��r�@��h�����Dc�������0��ɫG�_^&��Pv��ݻ"B��R|�B�F:�o�+q��e��O�\j:g�^��<[^�����/����'C�O���l�/v��Xs���%/�'%v�©� �啾�n��@y⑕ҷ;Nod$�ؒ[��{��Z"�
�X���3M��2>YG1�����#,+aR�ķ��]�P]�˅�����b�]E<Kwv��`�U}�폖�����]�ew�2s��̕i��+}�����A��E$=�P����������M)�Γ���xu�y�D�N�#8��͹�0�@�O;�ߣ_��V���$�A��+����*3혧�쵦�}8�'�W���_��9l���U]N����a�)*(�`����@+�����׍�} �@��M}�ͱ%
��S�����W��.N��4�1YB/��vP�N��[������ޠ+TqG��
f���谰fP�ll�n=^���4n�,/��	X`V
�e�{du�+��NsZ#F�>"gr0 %�&T��T`Ӥ5�|� �/���ϡ��/Q�r��Ή ��7=�Z)�}��.�C$�	��z ����-A����\mz|/z��{�9SZh*����Lڞ�q�iA��S���YH�H�b�!�a�IH#������Tp�09=�	�h@r0�=L]%nNbZL�#w���l�)�S����H޿ؒ��d���m@r�"hw�i�)�̋�2Yo��jk@�{`�������1<�L��l��$H�nT�vM\���y�My�Ie�@H0��Vҭ\�k'H�yOTF�#A�W22�խO���w�e��(9�Rn�@ꌧi���!=$��f"�7�@�!�5�4�8\��ԭ�a��f�f��ee1W�߭��>�܄Fo�q����|�TY�+�*"}d>��Fms��f�Oa��B�����%M�t~�ޭ���8Hkl:EM+
�+JÝq_M���d�-0"�M/�ؔj�[���VCb�h꥿�z)���l.�}��<�G�H޲}?�f;}�+�⥥s�W�y�h--�����ZF�(�~���?�n������Џ,"o?�Jk��,UZ�x��v��茍�U�N�k����s� -�Wօ��.;��Ӓ�J(TO�����n׈j7+Ò��o�;�`��h�5ګ|F��@ui�f"��lي��*����]��>��-��y�Wfq�㛆/�#*E���xN$f��d�����ׅ��
Jj���_gV�5ԕ���
��֕�땪�x��������b��i�)dyG����u���v>�Z��<!�)��_���Kߴ�����^��n;$%*^c�2B/���,=�����8Xq:][1����/��H=���:�|_M�����	r�b�4��"�����	(T�&N8p6&&�gE)\>��6���L�D����]���blC�y����g�A5�4�d���%0�2Z�Ӿ�ʪ(ڀ܁Iե���=�A$�u�5��	�M�}Q�d����NY������B�-���׻����X�j��a���)P��뿇�&)Eˑ�i��an���+�Mx9��tN�M�H'�0���WJ�9���vBt��!����u���6#,��G
�j�\�vm��@LU����r�sq��ߵ�;*�cb~K2�������9mgg7�������ű«�yLxKFW���ƞ�K~G\�dl�g���]\Ssa�3ɿ�ߨ��+p�LX��|�~���(���j�k��-�Y:i/Nz\O2��Х��}�7��V�.�����zX�3�LF-�^9�ir_������2�4�,�f�U�4�ǩ����ScI�i��y@����Q��NHvNN$�Ʀ�Q;��F
��6�b2/�,]}��O)|6�C��>���$"o;[.*�I���Q��4�t�b�q:d�&�PE
�Ν��(�<���2�nrfܾzu_�������	�J&�+G(7B���I l^>�{xG�r���"v�]��&?���v��U��S�J�+�X�^��d�Y��X���ȌQ��7�������[��Yvw�`}}:��,�v|�8R��ق�%[�h��:ٝF�_]�~6;y�١l���i{�N���A��޽
-َQ1�%7�8V80`r�R �nC�ve)_\��K>>��F�:��S�M��
y2���koW}J7$�<m����A^�ʥ��.����=�w��.+�bUC��}�I��f��� �`�8X,��hF&��h�#�������2U9G��YlK)���^�#RR��K�E���	/������1��/����r�7�>�EP��&�R7x@�p���ano/�s�xj�#CYF�t�f�zc�жc�*"�[�B�x	��1E�¶dIH2��Jn;_1]O�<�5W�C�=��G_�
d,{���Sڬ���-��mX�K޴iSI��0�n��{����
�TE�b|���"?��0�����|�	w�g�.�F#V��&�>��l'{�7[�]9m�Y ��%����[�6��Qr����,��2�DZ���\�����_<F=����y��۴�=(b��Vbx�F��[u�����H��\�c�=1�@{>�@_��aJ�'��!U��q8�al�ȑqz��W
s�v) J��9�=��~@Ѩ�~��N�p�v�)6�}T��f|'����`�*:��R25c��>2�&C��*za�`'$�̟�v�Ŭ�����A���.��,,�䣞�3�M|ؠ����	w[�W�}����
�B���a�"���`#�S��Ĭ�ج�;��£���0X�^�HiYq�ۄ�g�e�c�TI��
�4�M�+s�M���8IZϨ�PDr��ў�����K�w��d���Ҽ P�)%�\)���!��/**�^��}$�>/���G��;�l�v�˶SW�6�������D�w?�Ea�r"��u�K���v,e�HD�:E�tݤ���]Y�M��.�R�,�t��'�����n�|����^$e)N�E,�{��8���-_����;?-�4��߮�q�f��%��ڳa�%$Z�Flww���5H.1m��{�r��I�!l��;w���7�;���0L���O��k����9Ӟ��053#���<�)xLBb����:�) �)^��7���{��г���Ff��8&d�%�3݋Ǹ�n���$��I,���k�a�E��(��-X0��=�g�s@��8u.�����n-����z�Ny����� ��޹��G�AR�)e���r`�ᙃ��r�>J$������CO��B���~��Y�|3B�7'��t��1U�����54�pqq��� ���OOPaxA�t�ڳd^ }}�x�6�5�L��� �'&n�F�hfE
�� ����<��H���>5>&��hE���4���Uss����j�'�c̋�.0�ќ����L��B��;��<q�̈́q�d}0&B)��<h�ƍ���@�Ѫ���e��6�! #�w+&|�1J�9ި��/���Y!xF�X&(qp+P�,l������"bV�
I|h�)��ՍQ&A�e�V5�T�X�c-��f�g.�O�����F|�!!��@�xf��4�����Q��7�2��s,{��f�>�pbeeg�:������a������
��NzT���Z���x���@���-��2��}^���]�h󪲅��\�֡�1o�V@�7qq���uј$B1���d~��
~�F��y��#;[��x_|��j�hw��v�+Gl�Ϟ��k'@�� L_�a���.�I��)�l�w#Âa�c�O���8��-7X-�g.�BCp���nX8#{�9� ���HE�ջ�28!zޖF�{::\��+c�������h��ڪgnn�]E=ѹ<��S{�S!~�VLW�7��$�,��s�wtt�����\�c��{h4MVz�\�=s����6p�݇��===_à�����Փ��)���M4'��i%d�t�D�tyQ��d ���Ъ�<7�!�H��*�1D�6!M�d�ک����=@Y�e"|�#{����۱?�5��-���T�R���|��cf~aA�g�祀��y�> K�I��¾>&���#���jl�UE�h17O���vWtt�	3y���C����;x� V�H�G�Gr�����[G��J�op�m;�a�g��ҬR��=;����8��B#�@�c��1�o�n+�+҈u��7�b��8�SH�*k�WN�G�����d�q�����14Wֱ��lM�Vɢ��˄�S�a?�]����>�촶�����*)I�F�6��fؼ�4�hn��N���}�\+QT5��?�:�6��t�Tm�D�F>�v�3$d�m�V�fb��<1-M�gv����]��������JryW�:hh��x�UtG�?A�"���3����p�6��\h >ؒ��y7�j� %�)ioz���6�i��K���+�c��Qe|B!�bء����*����Փ��B�Wh�N����K�������'0ݍ�6��L��?N7m$P@�1&��%�'�FT�(��	:M�?��2���U���}�����k��� ?%����U�ꂉ�����������*TcҰ�R�/J�\��#pB�1U"*v'��T��H;~������-����0����=@}	��
ВA���>����=�F`rF���1�E�|(�SE��m�@����6�C�rtrR3vV
��|��sW�;lX�|�	_Aֈ]�3��i��?b���q!t/��[�����m�xs<�B@o������zu剷�� ��u?�Z�L��[����?E�����"f9f	�����A�8W5���>�jH�޼���y��h��OW����P{^��$�"�:����X�p�`Oqo\����`dQ�Ճ����C��6I-'�bd�-?T�e$���##����Kg�b�iy��چ���|.�!�m �ސ�wF���{DpP��q�%)��V^�́ժo��XҚ���:��.���w,�#A�<� ��9 G҈U
�G���8�0F�{d�i�6��J�0@^<�>�O�LA�# 6�����=�U��r�?��Z�?�`c*\�fFR��v�A%����� ���zК�;6��?.���ۢMS�(3c��%� �*��-F[�)���g�hy�f3��Խ�6}`x��/��:lO����Q/���n�w��bn2|��2�W�1��*�V&�Tَ4�Z&�SB�!x�{��E���b.\�t��r�;�%�N���m�����A�'T,��$hhG�=�y�hܔ�]��������rG�ٌh�_J���^����.���ܙ3�Z|�Fb՟ _>-`<�٘YY+:y�鍓�'_^0�j<h�H�[0{���~?m��7�g��I,ި���������I���n<5��1�����2�.ށ]��_�����
b�,^D�>tE��X�,�8����3�����Zئ�_jeq��4]ᤠ/��C0����2釉�;���V҆�R)�]� ���0)�d`�i?dsO2_������)E)�NI0w�%Q#]'�|�`�	��Yc�j���eה;�3I#���e$��r<���x�&KW)��Y�Wa�+��B	�;<+vF&B9�n��'ɽ���&���{ϕD/�����L()�hG�3;SE�RXx�WY�P��k�g �M���\(/	N�W@�`k�2xz�{�&���=	z{>{�Ī���x3]�DnS�5��4�VQ��R�m@ං،T�����4�`L�&���{���i{��S_��a�W/1�O�]�`o�w��Gц�ڒnj�+�D8HX��'f|�v�'jj��>p�5X�M��� ��|U]�B��K�6rG��b���F�0�#""\Y@�HU�����9�W2�\[��)���1�W�����梩f�ٙ��D��¨����m�)�����
�Qs��+n�זC2���������.?�aw�B�:����L��6,��w������x�VS�O�C���YԺ�=f���[00(�~Orr�2K����L��X��{�K�
���cOR�-����� * �֭�4�t\&�]�� ⛅O�
�ذx�4��f�(�߹uk-D��)���� 8x���͛K�*C$]�ª�u��}qNN�L*ku�\6�fJ�#��=(5����Z~���WBq�����/_qv���d�y4i�RD�Wp�c^�R[�T��U�q���ۏ�F��	Fb��ѣ�\gÊ ~������7.'�~~��3�1Ug� BQ�n�/�i�_`�9�O�I�[q�yR�~���H2tv��/��	�e(.��E�6�!���Pr�L���,���v��s�;]�b��z��0[�G՚��U��z�?=d��-#����\�2)2?�N���ÍIxM��s��son�[��a`�c�ð֧�2/�L�����7zA�Z?l�+H[�vv1U��۳m��W`�'o9v�ϝi1%0�k��F�b��zϟd�qzg�N҅�{aU���LR�`�`���7@��T���M����.��'D<yUR��o>�=�Em��?rL(�L4x~bo���(w�����6r�N���I�NEr�B��8m���<%��[��'��p�Iw�/Y'7P�%�������x�e����f��Sw�и������;��Mu����X����Ζ^�l���t�ȕ�����3ݎ����,��R��^GȪ��n݊�/`104�_��k2�Kx���8�n$%)|�Þ*���m-�"�zX�R����.�	�Ô�2��u]����v=!�`0������ß�c�l��,K��i����"�+��vc�I��\�4P�:3SϨ�ÞH�L,������"r:J�8_�Wd"tfEF>�L����� ����p�����$Yq����$V
�C���2 XՄ�)�t?)1���B�B�b��l?qq�7��V�>w1���n3O7�W��@x� 嶤-Ex�*��\������[&��7� xE�8D��G,�h~ZNP��M�SB����Y������� jO�QbN�e-���H������ `%��`��8��d�3$!����}*A��;@�G�l%\�.؄k�􉲜�<^?W(~�
�m.��<[�	��i|a�.S6nKӤ^�T!KכvڢQ��YM��a�y��/���$���������6r�b6�7f�Bv�'��í|����v��A�h�e��š��4֍nÌQ���K��G��,�Pc� ���ާ�Aߪ�����`>��q��"�Y�� $�ԩSy��||"�rHp��vb�@`�1-�����|����ĭݟ �xR;��c����^����;X]�����%��D��
�MF$mdl��~B�L>��&����&��0H�a�)<
���O�W��׫�5��*t�=? @��yk�E_���욨�+�q�uu~i/!��&�}K�`��m��ok���iʴ0*�΅����{�f��07��J��w7[�t�C?����,lYdAp�s��I�ֹM�F	�
,|����=������6���.�2���5y]�֮X��Tj&�d���*��:,�ȏ�9<����%u�.j�]�v�e����a�g��5m�N������jٖb��_�� ���:�2�=��@\"���g���KՔ��%��|}�fh�?FÂH��'\#'P��4IF��?Q��ٵK���<��)t��SXTTt��<��6[������2��a������ק�] SB����a��A.)z�9�p���Czk��X5���R�:����Ae�]���7p���
g��a^���C�����7�?�J���_��K]�W��G$��t�6ƪ��C���槭xpU�4�ʻ_g��ϱ./u�Hs�w�{M�����ux Q+��Ex
�2)�u	H8� S�
�t�/�7(_�����SkQ&8�Ç�Y�\+K�Sj��d9~u��\�q��VG�8ѕ��sr��ج����֔��\kJ B��
%�ӌħ��u��[�-MF>%v�y��^�ڗ�<?�4Bb�c�����aEz�Ios�t<:4-7�_lҮ����!��Mf�?��_;<Jp��R����x�w5��/��{� h0 �AJܙ�C�H�%����"�y��$� "�òt��FO�q����� �:��(�����<����]�W��>��.�LSK�,�|�o�����9�M� ��<��*g�N6Z��.���	����ծ�|�f�/�{�t�X��?��6»���Z�.�w���tϮ�.��Uu�����66�%� �Dn5�3��tU{�g�T�{2�D�E�2y��؅m��MN?u�����Q�U��<���c1{-�]]�!��t�zuz�U�<�5V�������R3NLL$M�"i˙!�ś��2K�� 9 v̆�u�r/�zI=H��u1��͕�0�т,���i�������b,�$*W��=�@� �O ���q�ͷ_�
�I�8o�z�VK�!�/М�S33���0�od&ӜMZ�AfھZ�G�lW�5��ķɥ;��V_"�v�͆��z�~ٹf�,�}#����ov�WZ�nd����a�������Ӊ/����������arP���,Tc l�tf����`�r�4ʋ��QO�ż��b���>H�6>->���C@j���,��e�}))�������o�myt��~�$dvq��^KP�L�'�ج�m�W��b�p�O���Y6��NҪ�-5���G��NM'����j�J��J{z���%6��r|�r[����f�����Aڡ�,���f�C|�y�w���/o����޼sl+�L�� *^�n���2��%K��)R#�4���2X6��֏�}9ߤ����+x�2.�abZ�,`@��4T/V���%]c(a��7<a�f�邚ȶ�S�XRK�QG��a(�3�MX�)S�č�:qi�
�����R�v�ik��rt5�*��'��v��aǘ�.�]�/ΑNL�C���:����[ Ɂ�sa������>а�5��0׈�/�*֫��M^|(\?QH�P�`����Ç���R&OA�cͰe�5G܁}�eD�C)�#6�o��`T����l�����y����@�!����x�ei�5��v�lW.����
���	WApG!�i֦v��������L�"���6��Q��ӳ?�-�Gn,22RE P͸�PӲ�eݲdH�K*"���c�����C�E�v ݸ; ��]�[��?�~�R���nA��OҴ� �q?"�thy�s�dn���E	iF�hrrz�2KM0:�@KeW�3���3LȚƋ����?.V�Bp�x�315WE���3r�\��c�/z�~>`F��ggٽ0��[��N`���S��P��ʂh��>��?ءw�(Z��h0���)Y�399�{^hrE�������%��"�������ץ����٬gGy����j���]Җ%&�	K��MCq�ef?F�c��_�빟<�4�����o�0!k��վ�2�7��2�s��`��?^�J5Vx��J�c��Y��lI ����	=�@��e��!���o>*C�<r��?�h�-Ja>r7ֱr��������S��vE�m�h��9w�)�{��]��_ʿ��߶la.׬��#�UbXG<_���d7�h[��y��7����$�rcQ�3���J�q�d��:8k��n�Fe�� o>Q1�HTR����z��ʪTzeeէ�Ƙ�߀_����b3H"�yg<	�N�%i�Ƶ����A
��lŚ�z�"ۑn��{����~��Ƃ�*1L�򆽎�h��YDx`��Y�^ܴy��#X����w�B����ğ��mt�R~�r�����+��y\����j-�#��oE�q�yze<�q�&��DJu�Ԙ��� &y�R�,f1x�4"��s���29vb-2u�ϗ�kע�'9�v�vt�]���G#v����4����	�;+�Ԟ"�_x��={��H�c�^��Xﾚ�D�ۀsC����>BySS�=5|7��Q7�R�����i@�'+ӳ.�g�-�BWE�ZѲ~�,�9�ng���=:\�2�;!3$k'ç��ꂠ9�Ֆ�硝�툛~~H��kݧr3f�u�8���^���jO�{-��o��v���@V���C�&d7���m�]����ɑ��Wó/����qi����W��d�nza>B+�e9��lm�bz@�;��o/*\����RO{� �*���"�y;�HY��t�I�mq��T"�K��t�,�:Zl�dd\�ZZ�@�:���콵��$t$X�_Cҫv[�$͝��@@��"���U��`������odM^(n�V|hx�j3�@E
���Z�IiF��U?l�{m�j<����+�~0s>&���q�R�yk����P'D����Wc��7~��⪅`I��ɧ�6��'NDG`��>���%NNe�8$`�x�$˗��� �Ng�ö���px�4GG�վh󪘪{�a�xyy9:���t�����^��O��_B] ��7��#|��B��˿�W���2-�����i�31�0s����T��(��u/p�`	3�G�[�Ҙ]����`/��o	:���	��Ǉ����rz=�N��N`n�P����j��x��\��ҵ{u�W\��މ/����v��� ITh���C��� �1[Y��)|xϞ����p?�J��d�G�n��&��mYV���7�8�B��l��4���T;0�����~�ؚ�Tx3lV(u�?4!����f����V����
?�=@���;u��e��ؑR���yٌ�kƶʍ9m8_a1�A�ѳ����s�� �Y���9ݤ��6�f�T�d������a1����Ax_�����^�i/ͻ��s��3���@`
f]�Y^���q3������s�~f�����8���ǹ^:��_k֮7is��sj�)�|�mq���Mw������ռ�}Z�@<1.��fz����i���^D�����R���rN�Ä<�[�M8��f@��_���d�� ��t��ޮ(�����_���_#R�O[?mgcS200�_p4�ʺ���m-)`���D����0̰3���i�F$�uUXn4pk�$3'}�	w�}���bڬ��rcmO�'{ܖ\��Fg� 5�X�P��?�l9�FUj�Ȟ1;=M*�Q��$:j�QUA����x,�mH�~�+ى���сr{'@%	*���	�zp X-@�8����C�nq���#Z�����C�R~�L:
��:W�ֱ5�����c�3�?��^A�1�v�x:��x�E�r���	F5��X�.�����8��'ؓ#F�qc+�'�" *� ��T��~�V�<f-'�:�7(]Y6qsv�Gs�N.ߠFq�`ǆ�y�6_	��c��9]�D�ښ��{�Z4��Ar\1����M��ã�6~��l]���uia��l4т����9�]v��=�ѕ�7�k�A��JQtJ���|ie�����l��ů�ܾP���D=^�D���,]o�dQ����)+��řV�?��[p�hZ���o���Kc�Q�@�}��Y��P�����FU
��h�2���xg.ʄ�p�R�� ���gNoA���+�����g[J��4rB?���X�Nf����Q��7vyɱ���,-����-�q���e��:������xX%q�;:XCfaayT��+x[zYĲ_��J���,c�t���1��]�(W��} ꖜ�Y60`�V�ø�:"�T��Q_H�o�N@�����iǡP�hX���X�Uk�AG�<���V\iC��+�kp���)+�z@ب���e�X�^yNN�!����[�WZ� �)s�ssW�e<W��&���,l �ucc�t��-ȭt�����U �.�g]w��e�Z%�G�l�IN"W{w���jQ�xL6*���P�|w��y,�~�L��Az���zÇ�lj'\��;v��m0&�%&&1
.�t0v�ZRE�]�䴶��6Ņ]llؒ��׀W��p�[a�=�l�y�Ȯ��X�|8}��@^�*�z��ږ��
sW�9a��̉I�����1!��%i���� �ϰ��1�4ܯ�V�h�����8��ݕ��Z�\$i�����a���缼pزߠ�<p�N��g��<pK��{��s���x����E[g3o�Azz�pS�
ox��\��[��Z���}5�w)�&���=���9������ޫ	x_�^�>Ӹ\��$��߻A؝�j�����k�I�Z�mڷp������]㛛{�������ݗ����;�R��~^���/����&�e��z��Go����(�Cڕ���4�d���+�m"�����B�Q��c^|���J��׻���BB�`�����ɰ񁮢�\��A�/�;v�<�å�������sp'{��%i�����tZt4������?8�Pe���>lQ��l�樯�M����&�?��'L�g��Nxz$��fUد��z�Å�A�q��ә]
 _i;��ׂb��r�&/O����g���K����9U[�j,8���Y?6�ћ���H�E�]s��=x��eJ�ȧjr�-AF��i��˯�s3Z��߹�ٿU��9��)w	a�-Z��ˉS֔�i��y��x���V�wG��G���b&=n���j*o�tPTT�Z���J�w<G�w�aL��s=�A����}�Z�2d����ǞkE�d�W}���_�ҡX�	E����t~�K����#���*akN^ay ��i��O՟����q���w�|�n�ڷ�3&?�p��3L�M?O_pD��ʥ�nJ&H�b�9J�ܥ;��'$�Zw<�}������c�~��s����Lѝ~o�����=���c;85X��Ln��d�o�a5�G̛�q`��`\�������ԥ84sڿ]>���汗Ns�]ͻL�U�/)Ӑ��1&_Y���}�(���#nǦ�=;�+�X�_�pџ�?��K����O��8���w�w>xI�v����I 5Xܟ�.N덜�b:{U/�o��9ⰵ?���>�{�A���9N=���B
L)�Ռ^3���wa��gnf�5(N��v���-O�s�x�=hI7�rf纏����W?j�0>������/e��-za:�b����{�k��������5ΘG��5ȍ��l�vy�V�7��1&�_���j\'P�����
;S?�m�k�gbb��4pu�{�����8u�FF\#bMk�Ӵ����7H�H���J��@���٤������`���|Ϟr?��̣�����-u���g8�K�D�]A��#v��_Ue���+��y8y�,�k��f��l������o9[2��%EWռ�7d�j���d�CSk��w�9̤�OoR�]���\dpD�C�tD�p	����_�s��I��kM�7lؐ�8�6��z��܇I)�G�v[F�O�2;�����*a����g��fh�!����p�'�r�˧W}�UH��>�rwE��cU���6?����0��qk݃+�Zo5�ut6HV��L�n�������Mo9�x���1��^��?dF��ҽ$ey�I�i~������G�!p����zS��)KO?��*��/c6��� {�y2F)LU$�Ar<7���� ������٤;����8��<=�����w��eFe���[�Ԩ���M߶�%K��(o����7}�?Wi����Y�����3�b��W�W�d��9mC_�UT+1�}*9�奤l���'1���Й���aw��g��x�x+h�5��uKD�nc��$��W+�z���K;N����r��
�g��A���D��-��k�v&q�m�-Uˈ-=�Ƨ泵�,cy����>x�-���~:���yzp:%{����gk	韖N�j+
��=��b#O��*��𒳡N\��w�4j+9"vҸ�=����uG��;"��/�V[['���	�&I����s��ǫ��6���`lM���zIQY�g�3�iv(�?��u��˻�i��.�R@���oUcM\\��9�������C�*:�����a�+��z�Z��G]���(�LO�tsVAd�id��L������)σΪ>���O�ˣ/��>����
�L�����=��e����ۼ�,3;�j� �?{Eo3S�p�F����7v����o�Iφ�-=����/������4ڜj��0�.�6�����R���p��}	z�jit��_��$ ����!Y�������`~P�m<�2c���8�$�k����x�n	Q��޼3YKA�Z� �����\�յ�~����t���<mӮ�<�9���7�x�ݹ�7^j�F����|Pz�9��{�ii�+��T���:��>���r����t�qю��M���A��בg|�s/p��!I�Y�G=~>>��'���&��g���Zh#��\�`LؽyE�VU	��SJ/�r�@k۬7���v���&''S�L�cZ¢������;�ͫ<�*˃�lb/�b"�1
�4�����=�I��= 䊨����,��ߨn�D_������p,����T�$IFG�
��le�gvvFh����l/�+�!!��MIVFF����}_�����s=׹N�����s>�w<F8DM�b���~<s�%��������Č쨳�S_S����"֓ٓD/����<7	��<����Q
m����hC�=�K�~\K� Q��7=e��{:����*-#�iA~���}F���hD~6Z����>��IG�:�������/�����b�2�ѽmQPD$�������@g�@�ӹI� [+Oi��L�� <��L�zg��S)ޫ�G��=��o�����ks��T����Mon�0{s���-���Or��h�X����:������r��N�_�
F�sTA�9^%���f�	�슌���zeBu����������{�K���oԉ�B��=��H�.O1F��`��Vj��~G��T_OQ����/�[(�NVp�b���+�MO�w�/<�Yj��C��Z�����b��ϓ��n�.r�"��"�_�$�IJb[����߅�����Ӑ(\��9�vs��P=����oԅ��F�B�kK�n��L�P]Q����>�}��R7�
JK �x��?=%/��V9p�'�q7z�ɉ D��Wo�{���B�}�6!1�B����)��|���)������mm7��4�Oy���5�T7��`?��8z�<T.^�(�}`>�m�sm�.^�"���_�!��gzĚo`b��־_��Z�������c����Vy�-)kG0�x��,��fa�#��	�iߕwB5~���^�Q��-�8����s��P���S�"��c���5���Nc˗��6���q�}�����pl����9�i�����n�����h�b�2~��'u�Lt���@�h��q��06��Y�H��R�zg&�*����)��1��)���	��o�OIVqfLN�%���v͛�{�g�����i>~���"�{��彩A�נB3��5���k?��sO����f �L�����I�����kP��U���������U� �Ag F��C�k�]���M��������s?�kfr@�:3_L��W�'�q�B���`T�@gg�6ɕ�J���G�D��3I�-^I}}�?�����
��jL�Ŀ|��#ÒjR�i��؜a����z����/7�gU�6��s�,�s*Y��Y�<��:E��W��P���{�����賓�����߬�!p�C$Q�nN�W�j��Y����aGʫ�ˣw����{��FMvq����Xx�E;!G�^A9�p�<�_�mp0�������''�B��|��!R�eN���}u��_	2�Z�p7Qx:1^t������f�&A���,q�ש4ҹta�%����p:����߮��<�
qz����bu퍊�D������Qξ���݇�޼��*��K����#��:$�O~{�ܽ�@��!�ԏ8hC�������{F��L���Ui��k6�rZ�7BЉOc˶|=e]��Cc�6/�D�H��{��s��S�vΏ��~*ė�*�����.����aA ��C|\��Q1|��9K�e
ܙ[�2<-[O������=�BK�����^*,g�;��;�`�����T��cK�<�Q���D1��t'vxH�߯��j6Zhw�`�6�-��P(���K��\?�.�����{�K��4<�Ć�,36�}6�����2'���y����������|q�}�&�ϼ�ӦW��Ry��lB���)�	��p�4I��/�c��g�M.���&k�(�?(N����isy���Ə"Zn!��{���:��Ӹ�����yj�P]`]r��O����$^B��+�A�C�,�iѨ�o�y9�$5L��#�	���zc���_��`�����_�ec��W/��1�`�>����$�`������:�
O^�SG���������f��L_�����f�4��H%v����/����D�|�F��k�89S��N�1��]5��:m��!w~6�_ ���q���2�MW]M9LxAQK���l�0G�J7Y�I�~]=��CJ���p�������Rm�D'YG��q�YT������6'7�!��f�Kh_T��]M��|{�o8����EMI
=�����_����_�4~?�@y�%lowp�c޸��S�F;���=�g���z����m�����w_k�jre �rӆ�̷KX�.�Mod�s�r'�� %ѻNb^���0\Z�.p������en�=AnR�lC<	߶���x��LJKο*!� 1#�U��M�cHW�9q~��qΔ����Զ͡��L�󝕄7U�'2N������Iݺ�"B��(�Hcؐ�cI�}�R\�C���f�{��t���
\�?��ü��;��P_��QL��X�{�ɵ��j�i D��,�[�/d��hO��9(���؟}(Â�?���uʸh����N�r��a�����'�����sE�ox�:�[��5��Kr���i;��;��;�)��w��G��	�~U{��9?�Sx��v-Ƿ*�p�+ �0!�1��묐?������]��ݿ�xl���G�|��bhl���Im��� :,�q���$���_�o�
��4ϝ;�,�9�O�0�JjN</|�^ۄ�\.��:�ȥY�B��h�L{�����1xE\.ؠ��k,c^�������V�7�^o�/���$�{��}�sR?�h��*�����Y�<��\��d�5֗����7S�>�ct������m#��W'P�p�����z���TI�"~$�C��~�3>|t"�6Y=U�nʈ�c�`�h����@j_��,���`\���X� ����c��qζ���'Z���6�A����d�6�o�=˶����&Pz�,Y�⟠�����P���Sh%*ɥ�Kr��[�xب,�J*̚�����������9h������v#�<�%B@�{��鹶	%�?yT4!%E���T�h�V� M�J8�>һs;3��I	י��鱵�t�]���ӿ�%��cup}}��Νݩ��_|�!w�����"sߌ�{����'t�8=�;�a����h@�)bzi��u5���J/yT��C��A��8�!G�Z&�*��<���7�Hdй���i������O�l�����'�ۯ���}�;y�Vi�M�b��fT@Eo�Mz�+�d]�v��d'��<��|�&�����W�v��W�Q�TU�{=W��<��ɦ͚9A"�X >����neg}_�{Z�]�'��e�0�#�^�r�#:>TS�co<(Uy�QP5�c;eX��,�B����=Ē��0	��P���9��Sd��_Zڨ(\�W~HR������K=�CRW'9g�(;ز�5���^*�[X�*h��Ə���lm$܍��ƅ����w��8��q*?I�bf#��
R6����ŕVT�XW>Oq5^I~=FA�v���CGnj�,��[���-���8
W�a^�F}/��z�MT�d��㕸�Z����OD�3����K�LF,N�9�
(t�o�'���Maˇ��-n�D�	�k�.�G�Ug_m`/>��v�)I:�$E�Qfއ;͆3�10ɝv���NZ&ݬb�QQ�i��i�d�S�{�	��&
'���ړX���@�J��U6��u:!�VYy1�����
���֥�q��|���o7�.�R���㶍�����p�T�St��Cn.����ȇ6���Ʉ����\��WJ� ��^�*)��e�����jGЕ�@��G�3N��{"��ݸ��ݟko>��|%�jw\��a26���l�7�s�J�6�]U(6Yi�:zݐ��/[ƺ�V��m��$�_P�NR�+���1$����~��8K}@��(���L�=�:Ÿ�FE��o��:��u��WD�B\�I�/1p�P��ipSnu��u#����Z�d�Fvj���ŵY�:�N�y�uG��|�j��=B>����$�mk��D��V�� ��[���4�;��'�h����#�� x����.̼��K�]U@#����vR*��.""R�RT�H]69%�5���$y`ʯ�����G%���^�/�7��rȰ��q҇�;99�:�^�e
�<{�ӱ5=��|T�%�p�`F*�ϩ��5�_�ܴu���!K�x��N�����L�Az�f	�n������_��o<d�&��[�y-�455˥qцN��>=��J&?�=���*>���+/+����-�3c��&�֪����s��E�v��l?3�k�PH׸o������(��c������z�C�$1ϩ�|�����2һ׼��{�4X�cu�A�ʜ�[v�:黎�mVn(��u40������H�uu�)㹄�� ��}.s�j�L���J-v{���ч����:y��os��-R��>ny�v͟>�*�U�ua�6G'7lYg���N��hP�]H�uU�v3�_	?���~L�k-zeU�A��ӽD�;3��"���	�*�	P\���x�pQ��f=��I=�mY����$qo��Ռ�̀��Y�n<���z�sdt"��dUԦbo��N�v�	^���&^o*6�ލ1�^�-����m_�����q�%-vzj?���j��ێ��IM13�_�u���s�-|uyhS������������F{8���Ƥ<�������=�?cވ>��yû�;m`m�u�qi�/���#Aq��kV����j��g\��7�ϱ��'2,GQ[gm����u�֓��2��x3�x2�ʆ���-�7n��AJ�%n�Qr&�ۑ������}/��Ctr<���K���/=E�V���?o�<�u���V���O�I����w�����E��ͼ���̕��=�� rvlل���蜦{6
�*_���]��ݳ�ؠ����I̸�����m$\8�~���&��e�Q�r�N�DҞp�-.u(�M�n��I�	��ڢ��`�ݜ�y�l$m��-�3�!�7ؿM�B�|vݎ��faeL����w/6���pr2.e7�۵������h쉼&sV5YH�b���X���K��#A������+b���;�(��!����n��Ι��:�7��&(�վ����%��îD����t��b�0)�t!�&mllB�k�g-����	�h;ym"=Τc}���{���bC��کjj�F:Ž�A�/��]b��Z�_պ족��D!'�s�U�L6�D��Pu���C��T
��d�K�/���:��������DH� ���5i't�f�4�
j�_�8_�L�9��Dr����L�b�~�'�z�)
���X�ʪ|���^�K����ָ52*��)	���0RڄN�ٻ
b�϶-��y����:���+N09m׌29�Pc����D���H�Wzhg�Wz�_�3�d%w���Ҫ!5��W���o����T�.�g�jRn[�PE�.t����iY���K^j�Ƅ7����s��� |岃��MTM��N�r\RU,�Bq
��IZ\����1ڪZ9.7J�R�J=�O>����這�C�4 �1���	�	�������:�Ie� �#�%�s�b�??�D(��h݌u�5(p��}���OYaQ��)
\5�'�0=�kd�1a:ame%.7��1�V(��Ԅ��P��j/���0eL��s$�Q�'x�@�|&-N������E�?ST� K�BKo��_��Q��ڐ����P����٭&A����{|(����5�m|�j6�'`X#�����>%V�CR��'�;��fAg@�p��t��ri�
�ͮ�^~���������IҒ���ȕzK�L@g�u��&;}���).|�ϑ�	%eeΨ�O��:;n���?%�2���,��&�m�)�7��R���D��"�}�4�QH/�"�p��+�x��6���}.��
&ٳ�������7L��Պq��i���˜@��$�g_�����L�M[GOq�	m�{����,4s���*Kb�o��/�(%�/-o����C/6�����ͪl��*�@7��dt���(���V��S�a�G^�Hlm.�Snm_������O 8f���[�����:ۿ��S��|��궷�b?D5��:�[�+�(���-��P�C���U��i��恱��E�~���Kl�)h���Ռ	��q��s�%?��R�2F�("�X�$����+�m�	 �+���L<:��uks}�xK���8�3���e/��ۅ|@WkS�i��Xp2$5[O+�����g�U{e�2��?���&3��)�I�h�du��]E^��'yau#��ln��he\S�#��<Ċf���7����'gʇuꆩ�;�57X�c��zM�,����:���V�S/ֆ��u�+Æ:���`�s̑=w�f¹�b 
���{�k�AH���	�4Y	
	�f_����<�vUa��'�����`
ϟ�O"�����Q0�v�6�� �8 �����u��*�!��ԝGQ�D�������.��Vsf���x�+,c����L�m�`��]Xm�]~���<��ْlP�S���T����EM(�j%r��9]Brr����/�#~9�{D8��U��0�*��l ���������I�JA�A.�YNql-�ې�������??\��i%pRr�W����"��PS�10�,9U�2�3�Z8���F���#,\�||ƼǾD.��N�ۃ��
>�ɹJ�J�pZ<\���(:�x�ȍ4�6�W���u4#^N�+2��.0�����\�-��+�l<E���$���c�ȇO|M��;�[RTD��\�ͽ��)�$
���t���O�K�c�Vs(���!���7π��7x���{��onڔ��46<��T]w¹��eEd�x���9Ӆ ��� ��yⓟ�����X����K^�ڼ�_���`q~x�r H���0�[���2�n*�|Մ�e�8c� Gm�Q��|ǃ&��Vd��w싱r��3>Q���}����͉<��9J��d?J�̛�A�,�ϔ/�����1�Ӛ.$#3s�'Y!�)�ZFb��2g���u�pa��ӛ������EW9��.�����.��v�e��K`�y2��}}}5�����T��7�W�HQ��j��@�3‧����i��� ����
~�����:��8���x�����9.VS<�~&|j����f��.�ȭ�L#޳�����$�ʮ�K�H� R��p ��we����Z����Rkgj6��O��~;��s$��,J�h����8J&���5滨��Y�§����]��Y�1�1�3����p鯿�Zq���KIu��^q��S��&�%�nLHH��>�?�ArQ�!R57�Q2���M��Pu��w='��x겇 ��a�������`��6� ��7d�ڄ���!��aZ�)u��jA�=��$$�'&�����@�&2mK��h�0��P��Hm��[�H9쵃��N�;e�ϡ����7k��`��!�r�w�D`�S�S��Ԟ�������a�d]����eLXYp��D��P����4L_�
 <÷:MJ��\v�nqE��1�Ǎ�ޒ�hfWb�	K䧝���t9�ʏnen�)��L�R' ��;����;�]Cè9���H��SKk9B�k��ݺ��|c쉰O�b,�ߝ��8�z�2����+�I�U{��M��\���)/S�ou6mU��:���¼�a��n-pR?�Sy�
GJ�Ebd��ZA��&R,�������Q��ĵ�/�
R�s����+ks)��/���:�?�Ҭ:^x3�S�<o�A�C��2��������{V�{�M-��4[����u_L9�qq7Ƒ3|�'m�`�2�}]賓%~�Xru	��>�9%�y* )A���������ǐ�1���]#)tk���>CU}���~�Q�x����b�5����2����3��o��5���J���g���ůt1Rt�,�l�1gᙳp��:u��?�)�[w e7�W����hjjB:(/�Q\���� 57�KjP�?�yb$��ai\q�r���̝(�<���� ������#Z�e���Mf�Oc�@���<��� ��ϕف�ԏ�l�R�(;?��k�۶�Q��!�b,'N��^�|m�?��S6���T�������b���0U'#�� �#�no����_�G��iUM�Zm��ˋ�9���VC��4u���i����lQב�����L^�Sg�k�V����լ,��m����E<p�E��e_ӺT:?=P��~m_B�L��W9�<is�+U�Z�<v�L��dʰӞ�q�c"���Zw��5P�w=�z����:�����w7	hF���~<D`�dChh�yc�S�4�N�(�u����,&��{�v��Ё��'�n�esi�8���� ��Q�|ß3q��$���a��B4�	 HG��O���ku��:^j��K�,��i���m�����AZ�����W�1�4�/e���6��S�|��}A*�6��ތMq�B�K�ē����z:>�l�d�"�zV幚T
�e1R��������l��S.���\ް(Q��k��X^^~=J����`�M���e�L�9���7�4�<�#G^[�Tm���y�w�K�0Ĭ!�Mԏ�C��t�:��~&����F���kN�W��,�{j�X�Bvz�=nO�^l�2O/���.��t9
�۲D>�9>�]�����hsH���%v��V�݌��-c�?h�}��h�
�B[��<�������c�AcA÷-jek��"�p=�A������64����V��|2s�A�s.�旑E��js붖nK��f��?�=Vȉ�C���)ᴸb:��J(�W�9��|Hh���4�!%�p��ʰ�B#-B*5����=�_�{qq��.{�H�����X�������/���5��%�������K�5֗��~H�խ�yl�-�3��>�a�H抃�C_O�~��ˠ��arP2A
3�V���@���&���:�K�x�����E_�_L�a�zU`�_F��+���8����k��5^�:���($�N]&����SI��� U�j�±�k��h��J!�66�Ї��M�	�8�} �O��ϟ���kg�i  0�_��n���l�˰�����k)۫̄�m��?���.�ޅ>s�a�E�M�co���**^3}B;�\�G
|~uZZZ���˛ߨ��͞�=�[��h�K*�N�qb~�����@Tᦣ���
�W�e#i�ND=��\c��GK��7�<ǚcΙzx3��'�hqY�A������Z\铓v'C\��3���9՝��%E�3��i��Z3[�#��-�;��D�&�|___,a1b�DB��\��u�~��T��d23E����9	Kn��c��%�N�n/��VU��k�Y�k��(Ґ`�%U,��)�鵅c���=��R�P �G4�;�۽�+�Y��[��~u���Ի�\;]��]��v��U%14����Ǩ�y��	b�뭭�ϖ2V�vd(�>2���.¸ۿ�J��UZ�ײ�@����C��)~��{.��g׽���sT�����UU0o�?��8�_�Z����UnQ�LNN�MǧO;&K&��/h�YWV6������E��Y��G�e�B$���zn���K���l�<o�CF�P;1�U����yK"���<�,�<Fd-E4�i� ��Y�j�� \ԏ>���ٱ��x��u{{��~��B&�{hԙJ��ȕ�ohU}� D��?t9o�Q6�rii>��r���/�qg��v�Ѝ5�������U$�b�Kf�|�(�x%���w�>66
�?��/�"�v�yϯ��de��2�е%��@���qr���$F5�1	z1[����e�]]���ʪ�����֜ԏ8�(��~� ���sysK����&SJ[�SYvv���]�x���s(�U�����?����n�Q��by�>5'�+��?aaa��9P���Z[[�R�8���V�6��CR$�_��tEKQ�S���`��e��A���s� 3���c��|@�/�QD7{�ױ�7�eL�ϯ�����E�{���`����ٙ�4��,�m�k+�}ܧƤ������dFƟ�����uy�min�SYd���4�͝��;�\�#�@9��W{�:`�zx�Wo1��վ{��Nx�M`K��0��z�uȚb��~;U�:��G����y�>�y�A�8P���ۋ�l��6Ŝ��G�� EEEe(̡��Qu��畼?ޕFu5�.Cm$f@KEb]��I��nC��/I�]���ᜉ�	��^��111`��ri �H7~�d���KY�:%������7IY��ĵ�$���9�Ž]Q
�Lz@��y��R���
��w�WDcZ�K�~kk��sR���T��(��2��WVZ�U�p�ޗ�0O�R����YJ�h@���oj���WR���YY�����)0���ͥw���S��a�sW��(�=Ĝĺ�+��:;9b���MV���瀨�)��������u�I8�I�s�֠4�ځ]����xJ��skj����0���Z�^@�o��;�"pl02x�-�gve-88gZ�f�~����/2�ɉ�\NLLLPH�Z���.6��i�M zK<-�:����s������Z����=�7R<F��A,���IO��a"CjL"��E�R)p�����#p�YB�j�}��{�h���!�G /X؈KU��vB���Av�9W�g��uujri4�����^GaH}x�&�����Ǐ�}�� ��G�C�A�xΪ���ru[U�l��'[3.�>]7\�Ǔ����u�>��������`��T������|�9	�{z��M'�N��\N�|E����%�1�'�)��f��/�Qx�tϔ`R���MĊ��w�~Lm�f�+5��CĊ�l��*�mi�S�e�I*X���r�8k}Y����p�p5��sݦ�O���M�%���|��+�}}�<���X��g�uPH�6�'�أ����g�w���y���o�Wh� �����|^�6�¡�������k�4'�$"�b�X���<������9�g�����]Z�=0�lR�^+A(%�,�]��_j�_�{�Ճ�j��~>>�h������*����AyF�ܺ�Z��u&���SQq�|�r���3$5���Y���3��n��� �������6b# ��1�G|w���� U��= دP�;��s�.�L��.��M���ʻo�(�Cg�� �T��L�yS��@�|�'�~7��`��Aon`��wȐ	@wM���ߒ0(s<Iذc$���.*ػ��Ƥ ������%�2�F��`�-	�A�~��j��3�������%u��[	H'��s�a�ڵ�f�9�,G��i����i����>�ַwpЄ2����X�a

B�댸Ujik�Ր�7p!� ���m�:?]�]
<\[k�ض[�����O���v�f�jVu�a��G��� �p[@Ʀ��aH�'�#�}H	*l��?�*�+RZ��9���-������ʱ��?o����YS�u @��z��j������A�h	:��*�[3�o7�(c\L�59��>|XV�A;���2p��2a���U�M���A�o&o<�.�pd?\��n��ek52��1B0��)��p������q�B�;�Vj�ف,��fe(P'Ooog��#��?W��ϟW�8�v�ߴ4⍃���(�|E��[���ְ N2���(>�?&a�f��Dt����Ç��zMJ��	#��oIpqsG��W���&cX�~��գĞ%�E�{
�A"zx|&��������cccP�_���]@k�1som���Vr��x㦋���kk�Nõƀ��H�f���#�`᪕!?P���%p�����8+�:�ekvv�h�Le��^�g�k��P.2�ձM���90�wΰ�"�Y"t\�Fy�w�����@�w��̴�p���h�^	�(�� :���f�&&�&������naq�X��N��/n:
.:
�5Ӟ-EZ��و���4_"�8Z��#�)����+��g��@�C�l]Z*<( �2F��e�/�{�N���q�*����7p��<m�t�D!�o54���k�wq!��YU=謭��Z $±c� �3�n���~p �M�:?�z�bY*�Mcf����rn�h	{���%j���89wv��5xh��W����y���������q��Ou�5g��!ii(��S���3��/�9�5�J#�/⣍��!�31u���>r�C��ݣ?yR�=�<��P�R���\�w) ��^(p�����2���9~���t�.Dc	^�щ!�=zgz0�8\3�v�Y��u*�����9A�}39�8�ר�Em�j�nnnNMOR��Y���mh�[U%���M[����kG��n�9hkU��`q^YI�#�%>�S�ҫ��Zr���
����g�D	�|���g�޷o�ǟ_��KKY����_�4�sRG��ۻ�����ghz9'?_�['����ܝ==Y�-��[8d���Y�?�X��Ç=㗑?����S�;~0���7��,�>����أ�:�L�2B=I*����ZO��������U��oy�2�Uɮ.�)�$��Ii��CKa��� �Ǿ����
rgsw)�"{:Y^]�s*ZL\\�9Ǐ+�І��6� ��0���G�}a�c+��˶���SSS�SCP��"`
v���ay<��!K$����fp��&JVb:ğ�B�B���Ag>)L�w���� �������'/�xH�4��Y(��便Bl�TK`�h��:��*��X�i�|FF3p�������q�|����*-��b�J��|} 'Q��號bd<�o��ȷ����]����;Q������i�!&h/:��Ǭ�J��ݞ&���:�Os��f�?!!��DDr�I0X7�$B<c���n鹼��%E��Q�AL�2��*�S��zϗ#�����:B�7��>Wɤ?u�s�U�e�7�����F��o�^^^^��yS�=}��ȋ��xZ������� ق��*I��yH`.=B���'�,�r���D{����ث��Ej|KK6}����Ȏ"몠X����0U�$ǌ��޶7��+�"&ְ<'#����K�������Ի�C����)�*t�D �h���9PM�ܪ3�va(���f*݃��7E���t�Vx6<��������;���j'�;�p8�m����ϐ�JSGL�򅱒t��U��NN1���4Kl�q����$I?HUnG$�Jؚ�x@�e��^�`��u��=`,�7�\��6?[��!�E������{���t��4`X ���!�<�NS�~uV��+��W��d��Q�̭�P��/����� kD�%?��ohٶ%k��F�$��kf������ཽ�s�TWn�E�A!!��o7��yf	��Ş�k���v��҄��3~>�Ga�,�DaD�U2q�j�b>���Ô�\��<�Natx�J�k�"�]]]�..��o�����":���~t��ڒHJ\!?91��*9tgUV�ࡀ�FE9��(����(���5��������H4`G�`�����C�[�h���X���a:EV��ϭ�-0��{����'��v�:�H��hiI�pcHJ��Ȗ�N.��Y�����Mԏ�O�q�n)*�_u���9��� ��0:�IM̌�#��F�����L�jռ�G�s��aSH����4�ݍi���@���o�.L=�����^ r4�����έ8,Ouӎj h�g��߿�]�a���rre)G{;;u&y�g�7�=��|
�n�ۛ�h��''�����V+I����?[�����$����Yp���Х&}q��;F�y* I0ߏ���d���Ǵw�.��c=�A����E��[�q=]CM�1K�A�߰����ʃ���Н׾�<]�:*�����a���J �	��'����y������9<(��FJ�6wK�����F?��]�S�-� �7X� 3F!�i��L�ݹt	#��w�''=PU����B��EK++�puH6PC�xL�km{\z�c��]/�#�]DY<3\g��gF���#���u����3?>�sEuZ����s��[[�E���Ԋ��0z�m�P��P��}��J������eX�������bԷY����,c���"Q}a	z�҈�1kB� r��M������A��� �6D Z��\�H�Uշ�04��?�ԦV�81�ʖ1of*�7S�M
t�fw.��_��)�el�mM������,�($j�	��Qƞ��ݭ��a��K��1A����kʘ�Z#�v�cd�WQ��O�"D���,
ʰ�BK(��&^m�f(�����v�c�/0v�����ۺ���g�ߑ̺�����|�7�09��]!��LPkOd�#j��D��	��A�*�/�9L�ǙX���A��/�3��)':�"g53�KKˏ-��F*�d����Ff��ؚkT�&��ֻh�D>��7����>��8���ȣ5[k�hyճ���6E� ��>�6(��ԑ犿�e��=5�3�9�����f���X�]IA���C0����_�@�A\����e-z	����/Q��� �|$����:��+W�i\ �uMok��k&E�=�7Q��ϋ5���`��i����~.��&��f�w����>�\E�Oz�z;�.�e&��V�j����oq��G5ѰWkz�cx��|v.�>��H��[�2O�ݽXk`-�*�� �֝�Nr1��!�'��?7(s�Gqk\��Is��CL{�1�x�a�Z���ZP�a�w�/���h�q��m��}qt���e�������j�`�p���+J�fDVm����p�n�	(�0�����ç��.b,ht.����7UPb��[�{Ṣ��䄺@�N}�-EJ������`�h�6�K�v�DV~~7��[�	@�ܤ !�+x���]�w���u�&K��@����ۅ��ۻ��8�r�@_��b�ȇ�	�i��nG(_mV�p@�߃��8���C��]Bc֔��%p��E�H��t%�_�e�AO��o�{N��P1�E/6iq�ߒȇ"�*��g��7&slQ}��R�#�� �E<�GHJ*�-�G�W�R��^G(?�C5~]CC_��1������+o.��u��6��ǀ�K{�����41�����:K$�X��M�� ����t������5&��d D�)��CA�P�����Ѧ1��8W����i�hU���ap�-�������|��]�or삂���W���v@��ywJ2�|�W�, �6����l������C�@h����c�n�����}���@��j�,����N'�)���{����Ԗ�Vj��
��<t$�Y��_��x������B���H@h���MQ����~���!�;��O�m���%��<_X�9�"�!F�zD?6��u4��S`�$F��F���(�fc����4�d�����h+�P�'EQ >���#�� ��A�P?�I��eU c�{.�.����#������B�^kq鴙��V�JKK[[.�B����S�l_3w{�1�ԉ�J!�P�t{�v_���0`ǨW=x{ep�1z�y�T������n?�����&h[�pXt] �h�I�$S�pKKK)<(['�{kO���/�)굹�-���";���d���2�~��~(#�3 �zP'�	h7�\\ 9�����ugT� >��Y̨�3��`҆lz��*2{
F�dU�ߛ��	�.���l�u��r��b��
@#��
����D�)����\k�H
��MF����u}hEjf�&�v�[�A�� ����E���0�=/'G�y��|��P�秈F���+M��s����ǏOe>��g�F{�� �e�F��(1��B-�|�\��!������!MU9��{{����������l�\7�|�+gaD�2ꐉT
�¥li'�<�2�6*�e	�-1��F�7N�ҁ ��qvg.B��J�aI�a%ǼX�1x;�m�7MF	�X$&ϝ;0-��6}p���!��X�q�-c�]/�؛���53��w�Y�T�h��s�\����U]@�:+���j�T�<�QM���9�����
��)m�j� ?�z�w	qR/�&��^���,��_�T��S�4�
�F!( ��6�9� �ޠ�@?��|2���P}��J$, �;/,�uV5��\�0�?qҭr�7�l�Rs�Jhf���n.U,���)����Iw������*M��������+uۛUc��
�����#�����_��Ä��Q����~���7*��p��%��7M��b���^�rJ..����H�������(�"�����ꘑ,-� p�U�f+�i2(WUs�����1f_��yxyM��&��Nr`:A$-��4j��a�Kp#�Z� n|e%p� x��8�{�s9jm*�s�!���7���y�H�q��HzUj��`�az�+�C���ZÄT6f�Ez�,��|�ׯfb1��.
C##/���@<�x�`Y�#µ$�$�_adc����ը�ӧ����j��lS�t�V��#�}46��ꦁ���3����(��E4���glчQ��%��IU!4mE�cS�[b�B;������%)�$wb���m.dT練IU�F��4�C�;Qxٞ��lm�(d���+��W,٣8�3�V-c�d@NqVT�^I��=��+F�x�|XlH�|�T�m���Kx���1��?�.xr��]@�*�$ IV{�r�3:�k�ϸ�~7�\5`!�_ -�z`����������S�&���O�F���+���c?wa\�m3!R�/����
jH6�ps�oxbD̀|��UUU��fz(F"#n��r/�N��!Cfac��>+����L�aG���/��U�a���Ч17r���(� �s�ږ?6h%���1)�?�1�U�WG)	+��+�����G�2��2q�[����m��
�1�q췿KQ�Ԍ#�s��~�� :� I�=�7���Y��2�7�.�9����d��p�7R��М�F��y��@�o\"�r7&�쓤��e9
���}������P�Wi��%����4�f�b;Hߵ	y�3� �Fh��GtF,����W�(v0��޹|:�z�}������188853��C�	!3��I��9@�y��;��IG�ST���[�����`%y�/Z,hZ��NM� ��~ q�s�u=�+�l��5 ?�9iiW���#hB���?tvuM���VQ��,<,<|jidBW�^�+�k���x%�*���Eg�3yB��9�]V��:+���䐆P�(L�ʻ�����ZTPD�i�fl����O��h\�pL ����{��ҁ�{�o�����e�Y;�3��L!�G���&_2�燆T�ˬ�`oN^jΡ�T��x��"�E��Ў�D@;��^���^�RK�TMD��àD��1o\		�b��ξ���h;���r^�Z	�D�A���I�L|}�
!nA���\��!ڛ�����[4��W� �K����A�L�n����m��<,]]]�#w�;;:,�1�@k�x��F��~�nD�Х�߷$�T�B��<ף��0@��k�g�*��+���M83��XF� �e#޸�w����JlZ靆�Zs�h<۹�Ś�R��HIؚ�(�5aɼ���%cE���!�U�%Y��h�{�p)[��B@ݰ�7�����jHH�S�B�c�%�4Hj��LN��Tf�7Œ���(=>�]b�c���zF�ӈ�E�3�Ä{*ʈ2t�-������H�4�z���Z�.W���ʰ�-Jo����&3�U�}�����%(�ă-�"��i�*́�\0�T����=EO_����8mF+&&��Ƽy-�|��.דQ�>tB�s"p����@4� �� ��c}�|zk}.��7~�r��VRQ��X]�����<h��Rmcn	���KK�K�*�1-c?7{0�*D�x�ҥ����]K�H��@7�@H$�/\G�	�ߛ������堼�?[@
?;$�Kz'�I�bCĪ���_�ҹ		����?@�9��q�D�B��Zً^bI��C��Z�����D�:NNX����y���0/fg���Q�����<��$2K6�y�Ə���N�����<~�?ʼ]���:A��mCx�|C(�S�/˙2�V	E��:�ќ�Z�L'@P:�u���)(�k���x� ��cn��!��&�UU����׫�S�R�/�{����'�k�Y� I�֙)ņ(0a8A�JH���a**#�ZY����$J���IEa�"Zx��XE[;���k� � �*���}3GV]����<�1��04[1J)�Oef��,*���EzffD�~jCb
�kN��/����u��� 4A&=|M"�!reW��59�a�:��hE[�3q�f�Yp��Q����������^SU�i���
m��b�DY	�2��8裷1h�֮�������H}���gO0�*�ٳ�PSR�;:���̱}��}��� ��`�;�\ �����wq��/ ,��^WW6PA-�,��O׉�R	;%�iv�
�4ik2a�<��k_x�I���EX�z���:z���+�ߒ��Ё��F�C�m�3jM7>uz�|������������|*�!�=0Ѩ�b�NOF�Fx�)�ٖs��[?T�U� x��Mc�/g\�'!�WOq鶕Z<�ScBL��
��vu4i��u��1�:Z��#�n]�e.��QҠs\��Sªe�0����G9`�3^đ�:���e;����%�To��c%�2�QR(�Ch�"�<��)�H�2��IHu��d�L�#!eH�B2d.Q���C��߿ǽO�:gkx׻�^{o��n~>��d ʮ��u�� �&�����`0����u6__�=B1�>��2\k����v�����p�@D:Gj�oŮ�گ��|(2�2��7߾=����'�"�e�A�I�K��@�Y�����`�qf�YY�Cʱ��i\~��&�_1o��Q�t������\��_����{䨪�<�QDx���ȿNnT ±L����6��?ξ��k�(:��^�j�Z�Z��H�~�9	�����9�~O $���}���š|7X��Fz����>'�yc�b>�)[�����]w����pt~�/��?�E��|��n]�n~QӏO&
�(w�C0<,Xq������\�"tk^9Gc��e]��{��B�/1�va���x�oh;�7L���ϯ�a�{qm=�3�Pm��`g�|� �2�8:�y��O��1��E�8�2���_s.����1�\ �~{�{������WRi-��;�O�� �*=,C/Ni;��j�y'��߽Gߜ�T�4X�� ����\��~����?ο�~~T�oq�o Xஞ?Z������l�-�]��Mk���6\�Yl���-�/`��¡��v"��z/�+���1^�u�!�r��	��3��(Zs��,�0�rL�=��-�j{��u6��y6Pd���f����$�g�C��J��>�+~�C~zE�i�w?�~��º�#G9o
(m	:�2=��ȥ��3����Ą��rS8��Eb�R�6��M/�_�_��і�Q���x�Q@�qq*+W��vÎ�1n�;#w�Uε���������r�^j��a�!�5��=З�dR�ҥQ��ĝ`��A
(���� ��I֊�.n�ԋt+r����[�XPH��+w� @��#~oU9�	���4���r=<,,�I�p����M��׿[_w��n�=�z��b��#u��#�m�_��f+/�	{.���ayG`mO�����&�e���U�M]����GTT0(m2���jd�H�,m=�R8��0�� ��|�9/�r�i��v��{��&#���a�^����c��=Ƶ�cƖ�%Me�l ��!�3e��5��SЊ���T�Q�\ �����Q��!��bCu��̻��¹�/l�����:���he2�2�x�7+�GQ,�����\��|ZȔ���_`���7���9�+�:r����ߖ�"�]����Q�yY����q##�OȽI+u�v~�6����G [�^x���X��p��-��m��{���z{<8�p��sO� ����������p����B1d, ��0�*@��ó_��f�@��4?�V�qz%IU͍���j�`oi94 &���D����RG��|1�X��.*�@/a1�m�D���eהk�$覴)����b^)[/�:���n��(�������#���
�Pz�Gutt4��6t��?���yS��&��2F���� ���ϟ?ҹI2��U���C*1�&?�/?��B_-n}t�-y9�,N+m���:Y��Zt�`��&x_Z�������P�U><\)���*������9B6<i���^XT��It�M�����`��G�_��{������s�]ʡ`��X�ƃ�ې��~6�6U���������v�����|b�tXm���h�6Mk뎴7i�e�1�_'s���������
�>^v!ݼ�av�!D�
H&�:?S��Ӄ4�OB�K��z�'H��]{����fF��+�Ph�z_�C�d]n2A�__��W�j{�h��8�"��r�o�����}A��3��Q��m�6l��7 �p�/��'�]�g�a�em���n���Y��{l��yI�0o�}��̸��&���o�kd�U�`����E�wYVF��b�g���싘��j�*߾�1�KdR�D0���e�_����:t��r*_��Ҽt���ކ,��o743���Դ�W����P��@���W��� L<��G�.�&'���	"�p(�?J0���@t�	d,�?��+Cr"|�a$�BƤ�8��ɚ�ˆ���p�ݗw��Y4jjk?{�����i�v��ޟ�x7y<�,�E�m�Y�O�6,�/y#˕=�Z���n�|�BB����.����ĉ�0Pp�-`6�:KB��7:�~<��ڟjQ������"}!�ئ�7T�5Y"���
	�M9�M扺 ^լaa�T��o8��M/،T��w���놆2�y'䖵��c&�,N&^��-W��M��*�q�+m|l`�u�ǏG�u��J066�����%d<��2;����nA�ϐ��ٔ�LF��#�ƪ�� ;��@,ܻ3�
��5x��K�`*�m�����4���32R�&|� W�t���܄D�6�g		���Y��#�4#�:]����lxvGv�����*��Pů�eN]j��/�~B�u(�����9�D�l6�khkG��jI[��x�L��f`]7�I.�����p~o�������6-��X>k�Һz/�8�YE�ӧ��c��4�͔2�<��]���ǚ�����~L4J��
�r�Hw�H���X[��q���T<�ܐ�Pfr|���(���{#cno�s��;&�n�wr�������*�z����N�AѵL;_�8�������Fr&o��Vsf�ǥ��_��ʲ��Ns���*�Bׅ�~]�/�tL�������d։���B�v�7AWrr�w�z�GeUՓ���@�jsv��p������l�H.�9j�j��t�=`����A�w �p�T�u��H6����p|����^z?���O�t�k_�Z*�:9��ɉ��5ww��9�ZL1�J;�
2�����艺o��z(��'_^� �p�4x�*������s~w��F�P��!�d:��G�M�����¯�]w�J��B01�����"1��&$�z�����6(�Ι~�S˛x4�(�������79�̴o��Pr�
��g�{�%�M��rĐ k/E�{�#\ggh�j�g�iQ7.��5��kn缩'@�|llL��`����"�@G�ɜW�Ź2���E&�MK�M��?��:�����A}�'~�;�I`��R������h;��{R���888t�?����^���ɱ�ɾ`�9jjiu���E,�������x|����rSM��Ǜ��k���e'K�P�L��y.�0^�U,P���j�U�����ɜ�Ef�N�v8+���n�[L��)+���p}�js�l�R�����C7zHQUՏS��)�����+B2�i��T$�� �=��UP���*��+
j-�Jz�v)�wl�������b��>�X��׮��ݵt�>�w}�a�9�5�)�1�eÆ}��K+ǆn�q���2��[2�&�#VC|۳�=t�Л���A����2j�j���6ۏ���]#�c�0)V�2|���Fp֔����,?'��ԏ����1ժ�~E5��Ɇ	��?�	4�2����}�`��T�|}}G��'�����(�'{!y���F��Z�j�,X O�O _��Eb���	Vk�D��8َ����1R���bd��e��w�T�ģ`XR������g�T�P�}$fQ��nk�@���j������h�		5�j��#���/�p���M<����Yk�yv��%R�n%�g���U���ޑ�����)��(���2|��]�T���T��ѭ��Ј��\B6䓊t�#1����[9!�c�&Mf���ڴ�IN��-<���t��󜤶J�l�xSW��u��k:t���V��F�K�n#1��߾}���s��#p��t��X�_��ű�~��:K��&.�S[�G�jq	���� p��T�v<������G]��k�l1�63��U�d��6^J�)&��b�הzQ?x�#���ֵ	Z {������3�f���D	II�H.J�K�5�?��*a^L=��!oN#7k	���M �p��,xeޒ�/N_�$�G3���iڴ����WQcc.n����������}�f���@��ޗ�'���{�]@��A��=���˛uɚ8�N�������K��`��|�B?�X,a�׸qe�-}��*��j�����)�	snY ����=�s���W�+�5c�P>4��[ׯ�r�W[]�{�#ŚF�����V,�8�[D*X��9H���ɡ�U�l�:�>���������������g��}ddd������
P���-x'�=	�`�CG���cV#������ݧA�:^ �e��`��K��5d�		)ӯ3<p�S�����g��;LZ��� Y]m6g�w�y��%���nZ�p�YCPx��� �����"��=�@&TƦ��G�eFD�{�y���Zy#���1��n4���=��Ku��F~�OƝ�9W�w��~qJ3-Z�î����/پ|�Y��	�Dq�����[�frVX��5��C�y��O���]����n_��v��]]]5<
&J��B^:���u��Z��$�L���|���{2N	�rh��ƲiP�R|a�"�����@ ��V�]��ȹ��R7:�?�a���ۛd}g|tT	�5��ԏՃ��ѵ�U����V$�g��`���4�
* V�y��3o������q�_B��whA�'<n��Ө��v��K&��#�*H,\M^��F���;{�g�$k��>\
�s㤢5�ߊ�5�{m����>��>�N�Ie9'��&��U)��E���#����3T��o��]Z��o�G��nDMH$.�9�?��i��2��\�p�H� ��y�y�*ס��5<�0�������1.��ц�@D�]�+�����6�����h��x>�F����O@Nl�Ui�4-X��3�^^�]�^GXL:�u���X)�4ɕ4��/|O)�O*H!���k�b��[#=��[H�}����emR~s���N�R���#���='w�.�'��4�w��D�����]"�����"y4>r(�k�����$��E\�		g�j���Y
������B����_��𥿽ie�WXX��yi=jB���Q�@����V	��9�� �l���0������'%���x��#��> ٳ�b�aӏ������u����8�<S-+��j������ey,�y|�k�f�!���\BB���`m���u��c�]- �C�ŧ(/]�x�cﬅ������-JR����a�=֗��j �;���Ѫ��n8�.u��ߥ�8TF�K]]B[��'���V��.���W��z+�}b�����B[���K��ן���KKK#.iij��^Y���P�5��OS�ֳ70��c	����ۮ`ۊ���Aaa��˱����{�V�M�5<s�A�z���_����t�O�������p)��;!<� V�P�<�'^?���%k��ȑ��uN��l	��V3����g�"�H��2Ӧ�6�U��C�?�v)�;�):R{6������X`\�4#���U&���&�8��s7Y��ϒ����Սq Nv�r	UF(�"6���h��>.[|�#��R7�b 0�K�ܼ���|1Xb��$99�y'/9��/xxP�~v���7��ߗ��_�!ر��� �^GȦ�/	�8'F@�7iD��h7����c����F�%V16��D?Ö:�ɇv��}��gz h!YYY�8�xr	��'Q��A0�81
���3�q��ڼ5ܷ^@��%��[�"�(^h �8W߹zI'=��d̩�$H�0����_p�ׯ_0l�7���m"��R��X�7xpX[Z"+��l��p���q����l��H��ƾ�Cy�쀛������27��wCI6��[��b$G;t�uyrŴ���&D��`��CDt��2���DF�_���`t� ��������IwVZ�QQ��u�^��AgXH�蛬�G�D�!w�n��������	��3����}��$���M��}����%��?K�0����w�Un��ԑ�.w�0�~<��̏�4��]	ET��cX���X`cҰ��(qXY9�v��#���g�%?#��� �a �n�÷����XƷ��� ��IE�MHa7����n<$-l�dݯ���/�:���DA���=����g;���Z�u��E&[���V'�8Sm�D˭�؁�`�NuC�������)���y;i��KǛmR(�6.�Z0Ȑ!���Ԕ�\Ν1�inum1b�Н� +w@S���~�`���С�����*f�o�_ ������ݳ�Ȃ9���<u�N�"�X�����'j�l�v� � D�3+��	��+H�(���kK�k'�Q<,�OS�&67FI3FJ��9�b	�|#~�Q���AT��e�B`�׀w��g���!�PH|������L]��뎬>˳v0w���.	���C��� |��0pi�b4\5߹���(hC;�RL�$'��9i���L���L�p�DP� 2�s'HK�gnB��Í㞆,���s�G����YDs�D�v<%Vq��+@;e��G�M鄼��""�\��g�X��=WX���i/^�H	ω�Cx��c�u=�:ܲ��q���h~O��m��XOJ_) r
[8�	ȰZ���_*lNe�jR`u����v���`���k���2Q.Cd01][[��U4S�p���X�h���i�w�$��t��UR�2�yP�#�l�F�r�yv g0��Y�mZ~b��j�����>��lf����F���j�C��2`N�[BU���G��.~�������5�D�E�ߗ�{�Ҭ�GJ���?���2�P��2	��{عO�29��J��K�.���r�+>y�R�&pA��Õ�h���o޼�O��
���ڪ�7m�'�����b5<��Q�}Q##��
��M��
�� E�X	�Nr���̑���&�y $S�����3�}<��˗�%GBw���ɂ!�K�����@���������'���7
�c[ed�pKi�ȏ}�;j���aR~���HC����i�Q4b~b�G�}+q�O��_]�S)�~�Y������֡7ϴb�jj�g���Ǔ��	�V������0� +�.H��s��0��l�J��<�;6Q����%n}L���~Uy��]�Њ�֛b�)>���.�7����V��j��$�22�$&��n��H��8@Ӵ�L]�hUjr��
6ρ/?�t������&�n�5!����m�c��_�׳��v=��߿���"�)���J�5iZlx%=}W�^J!)�
2M$}�M���E�+�����&dd� �0N��|��B��ӳ��,��/��iffV�C�Mț�:��:_�ĉG�E�%͢�C�g��ӗ%fER���p�3��G��Y��%���,�?Sx�"��`�f�փ?����ſM�CDV���`���0'Q�E�cz���㫿��T�hhh��i�.�K*���}M[������o;%����m��pVٸ���Q:70�¼Yl1����� ���g��c V�x��<o̴���i[��2B��C���Ϗz�V�$��OF��e�3�9w<	YS�=�2U����|�lJ=�y*�71�1~��72:��sr������ѩ�1t;��#s>���]�87���oV  w�!�+���(�f���Z�RF9xuﺶ�l^ o<p�ӑ�I`EK�qi��.7�,>E
��I�F!VB��{[��֋vE��d����5��x؁7:�.�x�0P7�Q��˗x�8�Ltٴ]���F�Oj�)E^�/�9׬Y�I���	�_���G���2���`R>~��~���y9��MC�3g���l6/�_�b��mp�	-#��}����OX�RQq�zb���?@��C�-P��4��:������iȬ ����M�r�[��b�-�F>4�%�@��&�v1�犾����Z>*������~�� X��=���)7�v���������n��o+�ș�^�Z_oM=qW���ǉ5�H�Uyt�-�IA�>�>B__�G}LK:5�̹M�! tOO_��ˌ=��eۻ����Eݥ
@��<��5�u��ub-�T	�B����x�=55<&
#�Rd1���
�i��JBN��0`[�͢^J.$]������(xCn��9�:̇�+D>i�ֵ�T)��y�Y{i:�y����ԅA/�V���I�K���d3�]}xs���C)�ׯ�|�soI�o }���� sC�+;�N�B�OO�� #������[@�h4��:����dރ�: }w�|�se �e��zhL���!���X�t�ҥm�� ��Ӭ���jj�D�����\^��Y~���L���Ԁ�H�8��ׄ�6 o�$i��Ջ��q�s����$9N6O���Ҷ�������������<����wG��ځ�� X޽6Z���Gÿ�|!�f�q���]Gbb�y��GU�4���Ŧȏ��wT|���~��� d��D�5A\�g��V�gu�����6��>%%%�E;33�Eܐ��?c��H{j�,�"c��ͧ��{鿅?�,>^KO/��4 ���S�!��].$��}&�KAwvԙF)ρ�K���Z<i��;�k��"4�����Aj9��X���k��sg��[�f�e=�O�EI�x��9#�x��F��۹��S���OLO�nkk��g�/���<�o`�D����Yk`�*⫴pה��~�Xё���ӬC�/�,;u/�� �gΗ������ƅ���%�&��a܄��@��w΁ �޽;\]S3&��x��A������MP+�o���:}�	 ��74�Lc��Ç�{a�sO�����i�����=��-W��t�}�(��!�ce%�37���\�WcX)�/��;26%-�4 >>P �T�rz�������x�!l�����Ss�˚��M_� �Ά0���Ξ?}� ��,6��i���U���NH���(�Wd�n��� �&iZh[��*�V�Ķ��ŋL��hoN�)	&#�2�k'Տ�7-���3K=>&���Ke��v��%�	�K:�[�bKEm�R���M���n�o�=����?>9�J��$�my�������iI�A������}e��
S��R�E�w�� �u����G}F9i�����"F6T��rhh(���wIH�� ����R��b�r�.�>S|��`�%�R(����݃37 �m[P	�ھ}W�'�z����P|{���F�OD�G ِ��HL�E�����p��8�$����Iv�)�3��H�,OǤ2����pIl����"a����C��N`\Dث�}}*`�M����;��׀�������������Íۍ����(I�!.G��hL	�`�QDI�m{G�Z$ԗ����9�ӴӦ>�����a�_k��R�@h`鎌��T�@�"0�������+^�)�潸Q�ބ!<OK_��d�]�O�N/y�h��O�t�O���ˊ}�K���q�΂��,"���=5#��k��U-���N���*GV~/���?s'sM�`ֱ��^���\�깐�׹�x50.�0Q~�3#�&���v�`:h7D@��Ǐ�.Z�$ X�0?�Y6���54.�i���V�^=gI�� �?}��|�x��*�w$&)y����=���###�E���v��<�v��6_E[����P�?AF�ٲ�a ���S��=HMo��E����]�B`A��f��u��=z��s�mii۟�F��T	<��1|���8;�XT�����HC���f�wgg�z�H��7,S�O?�^&�4�ge{�����/y�s��u��i�sg��^�L�#0�C#}�K �c�R~��e�"#�*����[��k�瀯!�R�A��Α�D`¨`C�7/�SE�|��W��(�����{&��<r���R9'}�����2-6�u�2�>\l�K���b#sY�� f�VF#^=o'�'H'�*�9��n�Ց���a�Ϸ?c�O�q��*�#S�������^F}���#h׺����K�g�P&CO�0�:r>�ii1qq%�Zb�����kJ3;uʲЇ|y% pPv<j:��
�f��m�ٗW�#X�a������ů��1m�SX��9̲9�Ep��*�]�:��<�Q'W��=7�pd$���;�DcHKK�	 VU|��sC�,�4T��Ĕy���P�X���f�Lu!���)y!��S��l���O��� �F� �� 	�Ωz8�����Ga��(
H��)��ɉ��4����E��T�Y�p���M�=�஌S�@k�v�'��̮�*�z����\�I�V��{a^��*�j�@qկ�<��U��<7��R��:	��%ȹf�Y����O�JH;p,���[G��r/t�?�Ek�|I	��S��ZSw4��'�{ׁg=��?��J����C��ҀSXO+�k��w��ie������0�u�%����OwW��$�2n�U与�Y�cl��KVU�­�}�����ѪT|�������E�����P�*X�dA�^�禔377ϖ�fX�>�~�L< T	*�!s��VP>.���jJ(��D�h*$ `ٍIj_���3�]��^YWW7w|'��v�B�)͗OF;������t kb�wn 1(-о��j|�����7�ֺ<��F�<�*�dFe2�GC蔊n���o\�(|z���0��L����I��wt�Da(���K���zD�~gC<�e���t�eй��C)%ϔkr;�e��`ֆ�'��O�fFm&E}��/�hg�p���[�<��,�����/$��0�xb����}9g𔨇�b��&�X�kC�r���n}S�ԿDLtai������kj����������RƘ��3�����9���P�}~���uS9Ӝ����h-c�(ط������
d>~���`�u^�6m:}�L�*�Ģ�;��3�����x�᠟��T�=>D_&�����jp�,0b�����ɏW��H$�&�<�/�j�6H?Hes|
qP�eͬsQ<4��9�R��K��;�j�#�����',��ڦO���(�ǎ��6]�k}
����]YYM�U���?6A��р�I��<
�]Fb�,���y�hO�q'����'/n���75����.�b��J�HB�a��8�}ۄFA����w�ϟ���N���9� v�]�1\�X��q�d���o{���|OO�±��S6? XM{��(U�3Ȁzěn÷�|Z� \Tf_��Aa��~��Ã`��Cŧ~���ߓv�2/��K��)�L�{��,!s��Y$�S�	j�1Ϟ�c��5��ꘄ�Ւ�Uߊ% �D�b�H�"}��#��A������� _�w���`ݾ�+�WlV9
#g[�0����O����ir��������s��s�!��0���yE����-C�8 Rn:,:S�
:���ӧO��|�x�1�}Hc�1�.վ �A!!�SChӁ�1��l�`o`0���RWD�ْ�>_,|a�q�=6�,&������D}N�(-qѵtk�|wA�����b��H\���Ш�u�m6��pnb��}�Ԥife�ڽ��G�z��-��t��b���ׯ��Ret$�#0�\�8�1I��z��PaZ�=̡Fό����x�YP@�	*�Z�{���P��|���|�w�ڋ����;�^rs�1/{*fq��u5V�
/b&#�c�=D�>&��2 4��(]p~�+Ȋ���K*k!X�,���A_a#B���޽{��ٽi�o,�Z!�y P�.lV�����d��ƅ����ץK/!��kP�4��-������E{v��$ǭ���t���h��\|��5~v�E�Ԟwj�K��K�����Y�VKHa�
kc�����C��P�/�����s��B�I��M��ÿt�ط*	��s�(���2NY���|r.wg��&Ar���s�IJ:�{���l�z���F�/4��<�y7s���ظ�S�>���TFc���? կ�B+Q
PzCZ$XN+p���_MuZ��`^FNN��Q��b�'��Y�yY��C��\��N�)���>�ym������;�T"ы�K�s��5�5��tp�D�/�X���N�\U���� ��a��@�ކ��[�</�\Tpr�Ԣ٫�F�%)�r" @�&ا@��s��=MMՄ�A�=v�׊���������}�����k�)�i�O�7|rjgq�k��@��R��&oo�̆:�˄�T�7����ƀ��c����]6w��-y���D��=x1|um��P��ġ��xf���	y���3u!���߂�0�z��ΰ��|J�w��4�'�ݕ� ��	��Ί��~2s��lć��
`��ҀI���<�|�_����&���\�|�1�K���)_�hx[��Y�V�*J���>��@��z�Cw[=�F����L��xtߑQ�����߿K s+��c߾��T�(���	n�~d�6��qL̡��x� �p��'�)���+_ZZ�UP��`_�(�$�Ű4��;\��2fyio�}�I	�������c��s�%�>�i޳kh�df�dfEu.8f���57�]G΁���U�1w����y�y�l<S76N,+S�a7ܜ�|h+�9=��x�O�8 FX �
�L��V�b<r�'q��)���>��^�"���� ��8���C'���O�뾸L+���QMh�����'��Sċ9�c1�l /�~����LPLLO@�W�]f�I���t��˗+���r�M3��=Q1l��:l;���` �X�2�A���3�#6��a��T�Wޫए�K�����;��-�o��� Г���p	<s(	UG�=�Ԣ�lܴ|A��u`����Kxf�ˬn)m��'�}��O/ߺm����k\�(�8��14�0`oh^����'��i
�>���z��B���w�p�pN�v�� �m<�>}���ns���#)�X�︊���=W�E�B�qW�Cc���L���N��;��|����lD�ٖ7X{g�	�IO�!1V56&�?��O�1�}������N�$]��r����:2~�������3�z%D?�B^'7:Y�k���� ��'b<��l��S�U#��q����@������EC��!#��C��'ΑU�*��ij�k�4�i=�8���bA��tڿJ�KZ��� ���MSȾ��9�H�RL�b	|����/���ȿf�^zo��]j[_�H�j����½]�q���N�'�2}�i6��c �rǁo�+)IU�׺Qp��3M_�k�y���̰�:v,���M-]ݧ�M�:�[�7:Q��!1�ͽ3� �½vVç�I����G%�����p���_�P>22R&��?��P|�)B82!���df�g�ͧ�Ok�%�~S�����)�|�����f�����>&�|Y[r�������C^������43sjǘm#���ϙƾ��OS��%9
 �⫪c4�����dUWV�_9�'���H�#�e���0':����y=��@IԦ+w���#�Ꜹ�FΛ;�����.~����� �VS]I���W�;S���591zo��7��J,���qjl��*E��9Q3ā�z�P�W��c��pU�L�x�=	嬬��!.$���X`V�����O�� u��)�z�\�#��E�@�1�GkZ�[tlG�, �<Р�M������]��ծ��Ճ�^���4��u�j%��
�z*sC�'����)=|c�!�]�~��%B��|�Y�zW��ĝq��p��[b}���EZ��˵����Wd���*c=cUF��w]�Lg��>~���<���MWel:	�`��S�l���`Π;w,���=q�)a� ������@X(7��#`�a��z����{��5�������t�]߯���+�q�c9�oii���,!1��7�
ֆϝ � ��RO Bifn�=l��x�ڢ�Qh'����6l��̭Ӛ=��G?�
�C
�s�����	Z�l|�������l�j�'0��K�cuM����;�Ұ��_iS4�cJ[��ǋhZ  j�U��d������M�0[q��TEO/75����XS�4��.R�gJ(DOo��������5��I��TjF4 l�ܹ�[��}�����k&-~��$�����I �)0�[�Np�Fn~^��G��_�~[X��\Fo�'y���{ϥ�T���թ���=�\֝��X�u���L��c��/k8Ԙo�$�tܽƉ��7k���ڞѬ�o�! ^�u������V�Q=��*�$����<<^999o��9��HAf);�����ʰ�&�3;pz���6ױ�"��x�.[f�ݯ��?0|l#�y��Ή1
!	��5]qn�iI�5�	��wc:��܆r�������D
��4,hd�5��%s�����l�5k�=z���Pw�	�ԛ�<Pq�5PM��Qs~8��H���&G��k=�V~��%k���Z�*jk�"""pN[8�b*��	��,/��t�p��Ȟ����p�5�uRΑ�$��� �1+L���(��}���W��i���;w.�40&%�R������V���/�x��T-��z4��}��W�h�`l�SO�Q�[j��}r���(GE�%K����⒒ѪBBk݆N�ʹH���AdR� �M�T�x2lm"�C�3�}b�yb�#�ի݊b��10"ҏl>y7ٜ��E��H,O�����~u�Z�5�<��,i)����5x�'�%������/��F«tAL�I��
.y`���-xuC�9����c���'��I�^�Y������z����w��?�c��,`�.�'�3t2{����Qk���p]� <5*㷆�?sVC$�w�^�����8��|����97{vvw{WTT覝�*�'!�XWKT4�L��eR7,=��/�X�f�*�	g��o�Y�8��r���-^-_'~|��tU�����h``��qWM���Fe*!�[*���}$�}j������|���S�gL���;�:B�DqH�_������Bϟ;�������Ñ�ݩ�X�/��_;q4%
S��̛���*���e�r�6���S*��Wnذ;|�������mt�Q%�$�f������[K�^������jM�8؍eY����	���sr�'��=�ÿ$;@%�!���]�}���t��v�n�H	�ft�-��ڧre�{d�Ђ7d(O�(V��Ek��c��ݴ·0�����7���@��������,��P���ɹ= �P�m��[���ÿڎih��.�;;6�!��8oi��tDޕ���]�%G��@؍��<�����*��o�!F�kǚ�����8l�OD���7tfzWӓ��&1w⢸�D��G}||�<�v���&��?9�CNN.�x^���������ud/x��r��&���N��:��t��.j;/��!s��IU8+feY)�-1�a�xkME}�j��Qѥ�{O�˭�wk���+g�\��O�t['�]����F���J���h�0���?_�U�] _
a�lr������v���G]Z���/�ǃt����m��&ɐ�����͠Q�
rs��<�P<]L���U��}h�|F��P
�+Dn�/�j�-�"?��(�����vq"w�;Rޱ�"����'Ё�}�~�Fy�OmY(��j��lrc����������I�u;��
�	G�
��FIػ�߾��V+Ry�!�j@=5=�]���]�V��<�!��D��HEc-K�m,s�0��fů�i��8�
&��߉��:���������ٺ�Ŵ��-�E���ƙ������W��d�+���8�_4m���<Ϙ�N�M�s����':��V�7��xr����C?�����y/8�o������Ԣ����@�bd'0�M���w�ΰ/^\���[�F�1tL{`�<	�C�-�`�R�'s~�#�������g��Ƿ�>79�[�;�>�Ym�R��%rw�[�~�N2R_�T�E���g�5���|IFfr L����^J�p�tG<����|�3�9:�}���u��Z���u�GF�ۀ�D/��| ��z�*��8�������|��h�&�D#�I��6���f�)��I���</�.�lE(-Zsi�v�!���iEc���{���@���� ���_o��^�y���+�d����r�W'ˆ�Z�[�b4b�� e�ޏWz9���HL���9�}Yפ{Wk�ހ"�Ы_oI�#����d�N��)��#$_[�Z�U?��i��1��,������ϯR��?���C-̟.m���%����x��s�T#fy4����kݸ���ϡ��bA����ɿ��&���֎T�C�n`�x�LQ�|= iM�?����/}n� �* �,������osfR�qп�5��Sq�I�GFG[�B�U�,K��q��	��L���L�Rt�<��0��.���J�po�QX�R}m��,D��L97��Q���|v�?6d2J� ��X=�r���d��5�t4��3�V�!h��X�SP�a!6���6�"Lf\B�.���n� ]|cq���o5���0
�iu����?�����A��<ΒK�½��	���\��+3!u�7����^0�-����s��A���߸��K��<�MYD=��@9�ļ>dz�3J�G�풓#1l.X~�p�p�~+�O�nW7�V���iI�2�	����$1+�WO���:3���-ɉ��ʐ�Ŭ (;[f$ɰ�gӯ¯�gct��5�t�̙�`Bc%�S��%��IXkc�>R��wf ��i�Mˣ���	��3-������6�d#��m�xӔ8�e���;,8�fz�.
�м2��9Mgr�^��n{�Gm�����?#k>�O�:X�ŻThsٌ�44-&TN5���?��孃@~pG��.���NL�����1�Y�qM~�m!��٘�ɷ�'��j���8�r:�X��N��-�m�8�6$te��*8�c��FAo�m����� ��0�6�XAw �?�?��؉���&�R�=�>h�cin�8	���>TU������9��C�2JvLq�t�m�BB��?���.���.�E�S������G�SI�0�L��o�1�?ZH엚^~P
�<���@�UZj*�@h�~��S�J.f"�^��Mw��N��5�����޸v�Z�?��@�o�8�5�8]�
@�N��2m.�Q�G��ZM�*�9%A��\ܐ�}d�1k���3�Xڡ�>(�R8[���%�	�u����V���:{�0�>�i~��a�;͙���������刍߶MM��@>�5H݂ �.t�"�����GsY �p�C.Ғ��t�^�M<�-�^�5.)����JD�"���|��
�[��L�3�m۫�*#�N6�	{'2==��^��2ߓIwILe7������y���`Fƴ�H��2*8:p�cF���Q�u�uLBB�Lt{o��8��F�X,�<s�L���bH�+*������~�.,X���}���OH��RQ ��U�s��)%��|�4E\�oC#Qm�k�;%�!օ����7�2�K�Ȉ.��6oR�M��8���Be J��dN}�FH<U������v[<}���^VB+��K��n��=߿�`�M�
�<��8�룋�ݳ�KXe���������*�Q��8u���kl����_/!V�yoA80*z�5�ʖKz��Y�g� q�hR=�����=�{cc��NvO�.�P��D�mZ�~�z��23�a�_�P�}�_2;����|�j7�#{&?d�>aaa�1�n���i�ijr-�8���!��;χ�ڐ��`�z��0Z�2A4���wV"Ȯ&N/����jz�$�
�L��&�M���眜������{bFL+�w�}���I��ro1(x���>�`��Q}��tEC���]�`dF�$(I�7�fJ�*Fjjj0�mF�R��*���zW�&4w%N7Tlkj
Q��Y�^���u}Dq�[���g9tDMk�-udd���ɽ��Aڂ'@+�b�t�F����ψ�l������қ\"�Tl�tT,�6�|�hu6Ǐ���; �@e�_��L���0X��zw�h��<�����+���M���c���] "�q�_H�de]ݪ���(�uK�O���.H9x�!��+�ٶz�� �F�������߿�  *FFn������ G��r����͞�?���l0+k٠B��X:-S�T��"|����D�=|�s�/v.;m.4���i8Ԉ�ݦhllL�hV�0���U����*�]ӟ*Z�Hջw�>�p9�������'����ʜ���b���9=0� @xA�ϟ� 5앥��sgZ�O����Q��d�{�R�VΛa$V��W���[b%�hق��B�W��9���iS�t�t�fP0õ'�"�;��A��z("��P�THj����7-`�T�ȝ�����-�M����߮�6w����/�K��8)1?&�˯US�<���\L��.�8�笀�r��g���}o�Vx�����!u�~�����L&�s!������h[�\�rl�Գ)0T	1{| ��>�aqέ��K����D���c���V}����!�!e���`�LN�.����w�]eZM��[j_�|���� ��@��ݻ�-]j�ċ��%o􊔼�n෯W==-{n{�L������*������/o����h C�TZ	tٴHX��J!��Ȣ�(d	�BNjZ�'''�6�웓�cim����677�ئ|�ĵ��7�OFc�>�Y�����8�t�>��D��<�Yjz�N���ģ�`�[!�E�K���>x��V����������@20��@�f��6��py^n��	���^��0�ǃ+0:\��o,\��ld�������t��.2�,-J"�#1�_��Ѳ���B�Y�ظ!zC�Y�B&���i��u�G%�\bH ?I.ÿp�̫%m��O}rA�qn�q��dkkH���00�6K:��_XЊ\~��[����n�;@Б`������o@+��s��n�A���&e�/����V��#���zմ���@}l'��K2ՀM��T�]h���O�N���d�v�a�" 
>�� <�M��]]^���0��ջl>5q.�r��-��-"B�q7����P#`����]�adOOߗ�S�&4�X�D?�����|M����>}�E�_FP��B�l8<�s���u ;��e�>q[�&����x�A=��"��í��o��ˡ�r�\Ļ|�s�mK���F0P�B��������bw�������mWˮ��7f?D�gF`X��*`��l�Rg���:x�D!�� nr��6�7�[�~���g����-y<�a3[0��n��>���Ba'k��e 	�.��\	����I c8���L��<g�i�b���zj2��́���2A�b�o��6NhR�޵?FDX̝��4-��)�MgO�?o�Ic���7���_��Jy����jժ�66��R�2N���v9�PyT"a.��k����\�����&�
�B�T2;�S���I�<ώS�Dʔ��$���n��3�e��3�w���������/g��s�^�Z�u?���¸�vsV��0]�jK�=�qp�p!�9�����\��$r����� ( a�{Q^��"�9J`Zg�WM1�UeeM
v��ia�Imu�A�� `�/
�X̢-�*�C9R2�>�2ӚW�-��r`3sss8��o�'���]B4Cv�^^�d
8~��OY�cT�)���y/� ����h��oݷ�>y�d/Á����J��-��X���MB�~�ԃ!����u�Rʏ�J[�d��OP����)���6�*�i:���|^�Ao�|�c�Y���ӎW�<�ry�-e�Hi	�ŔNH*6t��;���A I��>\�'��Lu�&�@^���-�����wu�u�I�a#W@-��34�wY�ms-.�6�nhbT�jaT!w�3�1�,IZJǡG��:�Z�v�a�Q��k;�I*�O#S�Xhw% ���4�CSwc�Xx�i��x(\���Ҳ�j��ȹ^1���
�5,,����w@�9���1�8�%!!KΥ��j�Fr
-q�%�����!�:�_�F�W��)Sdɢo�9�������e�e�s	|��W��k����,�� ��̀	d�$t}��5��]Gk�����D�x���|Ȉ#w+�'�!++�OmP��ò�%����16�\�Wu����R���S9����0��Z;(����y|ͪfa�Yp#���\˹~�$ƗqdM:zzy�ڄ��WS����7cjkϓ��Xr��� 3u����G}�Ʈ�Q��x��ִ�tͅ��=����l���~�@�Lk1U|����GC� <��.-=�e˂���?e``��(ר���]�lvB6ݼߕ�M����rճD�q��jvߑ��!�7��(��T������ݳ8+I����	qꍖ={�����ft���*�qqq�x1$���8��r��EY��+��`{��:�:�q��&^Im������7���-.,���@+z��������t�+[�J�$��a���'wRT�BU�x�:.·w�&�S>�Ҥ�˷��kt�Y��N1㗅�/*�����K���9�g�����\c��Q�eEL�����M�g/0L�#I @�B��!j�OIr�Ww�������M���N��^
�#����h������I7�/��|r��w�L�<A�*~~
�YB^�͐��/G]�6�^�b�l7��ހ��&k/��Vn���b�uh\m0��4D)eO����[��&o�hyww���Rn4e�UW��xU���x�w��ˑ�%!E�G�� 0�`h��Z��XA�A�".�N�Yʓ��k8�tB���餴�a�s/眡9 ^0~��w�_�6��3F7+S���zr?�)���⓾�l�<A\��ek��g��Ţ�����Fm�]��0V���+����ԥ�5������gl3����HW��;7��9�). ���/�E|�);�f��#WUU�_Us�^���H�E�i=�n޺�T�IyM�r�����[�eg3::�����I�㫸!��%ෟ�(���"\���P�,���bZcT'�Ny� 0�8����7����O����Ʌ�,5�(���!`��ٳȶ����&*	R���ױu66�=��q���%�]�aE��a ��7�Nn�~��l��^p�]滇�b\��R��Fݥa���m��\w'���$/�} /�H�1ta���ج�f��O^l�5�|�^l�YS�\ t����@�cR;�Aoˠ��T�:ʚ�1O����--O,�����q�C����ݔ�S����SP����"q����a����~�F����TUV�ƒ��o� [��i�[@Bnpὥ�]��2�����X&Ld)S����,��/�5jи�+���Sa��--���\��qǉh!?���C�D��C�Qv�r��7��{M�[����7����.��s�n�̱jԨh��?���Aު�7t��3&���w�#� P蔶G"��@� �a�v\����_�(��"ۦ��>7g��аPW`�U-�`�]ܖ�R��"OKؽ�yX�.���L�w��z�|���o)F������5��-5�EFզ?qq�f���<1������ |b&����GiC���W q���
q������Y:�~?nk���hB�235���4�EȺ����0.��o���`@�}��$��quu��y� u�d�P0lѩ���'�1;�*r{�ې��w{z»x6��J8�����B����(TmC�	+$���I�ס����� 5�a^o@4z������5333����yy�p�3�zAƅ����d͏?��&���O��3�Z�G�[�Y��k\�-��Zs�Z�N���,)'k�b�Rz�毄�dPu��ٓ�
�8�"bA��$��	�>�%��i'CC��C��ۉ��� �DA�^�elll�+4΢}���' xV]A��j$���b��)u��-4#
�%���^s���U���*�5�E�j�7��fh;#�Τ۵ ю�)��m�=K^���-�h،����(�j�}����-�B���k�T�\�y���^�~�ݘ�m�O��!���2V��G�#�����W�I�M�B�d�+��E�p�M�.���^W�3~��n��D��dj���?:
M�Țȼ��Pʰ4j���_^.C�ۈpxP5�(� ��f�f;��.�d��SVV-=�	>� �H�@��W�7��D��:�4;9�6�󤘘�<"֢�Z�#�"{�����	���f�\�HY!I����������y� �,dl��
�@7i/-�,W���?&��pp�Ɓ([ �-;�w���d烇X�`�e}����P.�6�$�����.BJ�CI��@࿦"�-$GV���5*K���͚l��ic��_8;5��D�~��D!�=kћr���O�Nۑ"\�����7�����GmB�w�G���P�^��*�(��,۷C��GE[$	,��i���Ve� 	0j;�r������5���``N�0� ႁ�<�Z����D�N�iB�p�%�R�^;;�Hy�[��'7�SfV�҇�yڨ�*!UNQ�y�Ĭ�3hܳ�ewvv�@�nyz�y��/�y, Yʏ�t��n��
�����@\^C�Ӌu?pB���ID!;����܍������b�h�3;�l},�����F��Ƃ�'����(����BhZD��A���D��ᖁ����^��A�w7��mも8GCk�Z�g�q�^PXD����Ӣ��,v�����G�!Qÿ�t+�zv �sݸ^BRtS��.B�H\��+�L8s��a%W)��I!O�0����$ ����=Z�E�u>���9ȢI�aq_lEhl,�e���l02)�}.쯿�"�\yBE���3�H��ʲ>n�0�a^(�ښ�h�̶�R<�1�v*�.�#E`�
�9'׋1Q�p� Ty+����Y���Ť?�Mc|��ڊs�Д�ɔ�ag!�S Ehs��� �	�����ؼ9"*�S������CD����m&�g��Ͱnjg�^����6���yӄ���ڹ�&]%}��O�HJP��W�������:��[��]�*��p�^��a��B��U��'=�k�^^KVڹz�L��>N�s�R�:$3-qf�a����ؚ����
l8��t��$�~�4n&x�̸����������;�HJn�d�����_�˫��O���653�DK��B�	y��͛n�PfoμW�1�d]�L�{������U�zzhi�b���|cpA��7�O-1 ���/υ�7~eQ�KJ�L��A.x/p*ـ��o�k:fAL�'�����d>az���_��
p�4&�L����׍�࠱��.��S]�A��J^6��P�]��4����~���YBY���˗!{B������A0�|k�<��Md��틻�!�i��	a2�[�����K��K��j�s�!�F�3yS�@�[:��y��9{ԯ��Bl��7멐�l3�B��_�>ыI��W[�j҅�F������,6���4i֕�oa�e�s��Z�����օ����ߵ^|RS��E��8�o=�ɵ�&�lVW_�%�SJ�����%�CVRJ�3�.a�j ����)�������	�� eO	����.[L�S,B�Z�9��>݃,�5����ӳ�F�lS�9�/����ޛ
�k`p����t��i�	~|�ۓ���(�J
/[Ԛ����P �<� �ŁB�DO9�U��׃«�Yy�{v�G�r?�K�ý!>��� [t�|���( �-"##�{�F�a�h/*a��Gi77�pj�o�/����Cv���>����������;����S�����k��D�����`��e�4x�y!��3�����Pг�v�_��D|$rr����4�ir�HS������;uOI$��'��č{N��g��v-ҷ�
���fgvJ�l��f;�t�G{�ns[y�:l��+�&�~Z���~�:�����ނ:��إ��D��"�wڜ\AcM�VT���o�� {tK�?ioH5$�p�����{K#�&�X�������fo 6�Á!�9�����t7���W=��+"�^�����p�1�����	e�[`�~!�5�߸'�vm�a��;Ӈ��Nn��#e͐�\ٺt�֨����_B�ۏ�>ccc���{���W���b�#AP9|����4�?����٥Pg��)�d s�g�"���v�>��M�o|�����/>>�v�"�8B|�Kym��*K
�j�)~�;L$�<:0e�󬰰���x{U1.,`^)&�����1�>Pboo�-y$������Ե� ��<���(���s~� tZ]�ABF�C_����O}d��,{!�\6�����!�]�^f5j�,:�������H0��"�wKE�,��wo=G0�����F�[��+/>F~9?B�PPP`�i��0�֭�?at6&&��޽{��D�� ���؃��F����|��w�D�����S�4���4s;��g�����_dU�:�1Vp����D�3r�/E>U6�<6ߪ>�!��a'�+�U���T�&� ����Y@@Ey9��0�|����� ?Sè�)�b�}2�6�"�o�q�b�~� ^Qm\q^0\������n�=��p����T�5MM����A����<<&�l�^[[�Lh	�o{wP9�`WIH	�`n��f��x?ga�`l7��c�!��+(��R�A<���Fq�Q�`pk���OL�n��r�x���uȫxf�جg�O֪�qH���l"IP!�ߐ��,�~�T'vAgvrH)^Kz��ا��HY\��Kb~
R�����O5��^B`����=�|)b��è�T������&�4?
���%,H����/E�����)y2+����x����D,u�3@^M�L^�0�=R�
�;
L���'���oH��Q�o�q�@�sI0�����n��r��&�	��@�0Q���4Y������xw��9�/R>b���3��_<�=��HoTl'�N[x9u�<#p������>Aj�N��_�S@��W���v���<�����D�^��
�1�_b�?���$텪�Rg��b�� ����!��=>�UңL�LO�Q���_6XEk3�J�V�����&&&�����oU��cV-N��cU�?�a0\�Gyno&�!o���czv˝�A4Z`s�Y��旇�ώE}ݯ�F'N?��K,�%I����Z�C?�qx��R6npݕO�F�W����?jѼ�
��8��e` ʄ�;�~$�dAU`���l��>�,P%м������׽W�S#�$���H[����羢@���|N`���`CJ��y������U��V��U�t[��y�c�pT�Ƥ��D,��غ�С$��Eqd �Ԗ�D\��޺�)��v�lllf��D��6��a�����VC�嫄K���v��X���3�Px�Y,H� �U��⩥3�@�i��"Yd i@D1���G��w =s��
ѣ{�]�jR?�J@r�]�Kl�U}��m(b�s|��XlG_p���駿Y��5�l��]�3���oZ��'�4:�@y�Pk�<��i=֓��xwŧq�����%�JĎ�Y��X��G���3�r��J��.��/ y��B2>Q���v���p
���:��S�_lH�οU�&��N��fVo`���n�ϫW�p},$|�tSiIUMM�Z�ɿ�����.]4
�.�;���+P�!L�A���B�C>"���R��h��q�P'�}[�	MR����Y�� ���>x)�Č��At��Kn!�q������5�G@����p|ρ\C�1����,���;�531�0C����p�0��fL)�8'%%e>Ф
=Z��#�^� �	�g-��T.�{�����d-�D�"�2 �lOY��"�0v�������d��h�]�iRn�9��k��\�&L�y�?���f
�\����ʪ���Uʹm�v����vN�<yY1oJ�v����-T�h�VJ��%h��ޞ�޴A�c"2��%7�+���ӊ����ۯ�=	�6)d��c��&��"�B�����#�T��ROT40�222����/{;˒��gjKn4�A���|�͠�M�Z�jk�qE�G���� 0��=y��jbLMM��^/���1�|6����!~RA��xG��Dnh
��(�@x�TZVSS2���[}rW����aFډ� �%�l^{�6EPI�F�'�H~؉�PJL���o�h���|�8	����sD�,� i�6gcc�)���P$�P��I�yMڹj�̧����|�f^J?9�sE9A���`�@O����o�>��yyx�b��b�7���m۶�o���f&��&p�U����O�O�4�)�@�����d3!�@@����4�t!��jT}���p6�
�Q���$
��OdC�F�`�e� �>?9"��)���
�7�yTP+ ��V����n} �G��Bŭ�1=Y֙`]����.,l�Y#h��s�QMooo�Tcmԥ�Lđ�6�al�Yq)�� �`^�P�?FR����^?�PZQ�Ѷ���}�.�rU�!S�o�,��|
dW}�em�����q��H����ʤ��V���
��y�" c�p������3\[b<d�2�A�ݾ�8M)����>���K25���-�+��,�;��؅����T�8cc�;?����~q8��\�x���Sȴ[�LZr=JB��.tv��ܔ�}���E|�S��H����f�ׅTVW����Z��[�6i!���ë��p�B��.���鯯/���j=z�����R6�w��Hun���\�=��X�
V�폌�.p�6�b��R���c��7LSi��	�dJ�Y�|�/>]��p���SD$ip�W��I=ڑ7Ԗ�vao9��q��dd8�1<<<�QRb��c�Dtt43y�Sٜ�;/d��9�@E"6f <���s��m�st��O�w�����	2��V.���� K�mO�7�56k��<����W��!Q\�E������L�w��	�����#�.�h�b��8�!>�'ۉ�Ɨ��n�����3 Ԏ� �@� g1s��\�>�>?�=/�n��-�z��'s�w��&]����R�I� Q{w:��@@b�X����i�jbe�tK𚇡֜�o��><��K�C�-89q>�x�c)v�������<�O��o(�H2�*B�:��hW�JG"z
�rqad˯���
��8��g����$�FGl8�h��R�$�F����y��ā<r�!�0 ?x�j�z a�o����@��c��F�<��OVS�#�%Z#�EPK�\L�t/V�����#���ő}�3�qf����C"O �	����5 �WJ�u�J���D@I���t�D��a��y�S�Ne{Ǿ��!нʴ���)�K�I��G9zo��W�-<�]�/yK7��{֋�)	>~vWȤ����Uk/q{77u�JjL�r w�L�06<i�@�Q.��K�Uf�_�t���+'��Sa8�e�\⃮z�]D��g5^�3�y�l��8�S]DǑN�6�t�@����^�k0c�3�i��#^������O��N4�X�R�f7��@��Px���VEA\#"�{lԧ -hP�UsM��l��mhr,p}���,��=�>�N���'9��(��$dV�ӫn�aV?��_װ��v�7�.4/$�����	�~R3~mV��UĎ��ԨUG���d�2ż��>,=]D���en���92�4�GP�����mO�۷?�E?ĂlSN�/zvLo�O}^S�zH-��8G�����Y4����q��.+6�0�_�h���
@���c���H�A�Y��!6���"��HM��&�~"�s
�� -j3�LԬ{�q˻����Ǯ�@�0\�Ϡ�����!ߛ'h�QAA���*�d� �F�#8+�y)���NN�o���� �I7h���Xz��V�Aќ���fͅ'}\�zյX��& �Z^�/vٺ
R�e��\����`�NT��zl;|�o�	��t����K'�7�S7
��ޜq��0�/���i2@لX�*� `c~S�M0(�K���x9`i��
`,��X�\]�>��Ԯ�����m@"}��F�JJ@
8�gq�1h%��?�(�ع"��i'�ֳ]�!�?�W;��%h���^t`� ��1�],�����qJ	r�����H�>_� ��<t���_��͋( '���y��=W�����!�m)�y!�y!Z@K���9���g�l�
�C�I�5j#F�9��q!pK����f�t�sF,PK<����]f��yr2s�Jf�U~����m�S�L��o�+j�=���d��ma�	��ܞB��B����z��^�%]PP��usyMӎ�%����vf��APǖ��s�|߂�C��x��=��t@O��:�kY��)L�0�x	���o�fpQ�����}.k�U���D(pg�THB�'4�T��-����� �q��6�w����)-V^�W"��|�1������x/C��	r4`�����^�\�wI̺���von�<���6"�	��ː^@f�N��`p�bQQ�UbM�f�#<W��,oNw����s�AF(~��p	��ϑ����;u�N��^�u% U#�|:]�A��m��!0'=~�U\\�5g�^�10��� O�k����P�^���1ș~�H���X4���Z��5۹n�*Uh��Y�e�c^�QJ���{��RǪ�M��F���WG+WTW_1e��I�������q+R5%�I�s�Y%V#ͅ��K���Grc���ZGr(@'2/�Б:�X\�[�����M���8�%DN� ������9��O�AD�W�*�j��vs�XWI���=ni2�,���������|��a�@䍍�����L\���<��J8�= �:r��@��?������3����1����z�������,[^GF�M��.��5�G��������v�k1�C/]���ZgkApiiF�����W�g$�<�K��8�E��X��\�t�~�Q��):0�8��'��H�~��#�]vX�S6�����\����/���逵��b�&^�sL���2��!4�cѢ'�h;0�^]����x�I2�cйZ�o��O�S�Ĭv��!V���m	�}0�g�����^�*�@f�A)"�~����X�6]]]��w��M:ρ6Y3)bi~��.�[�wcmt����E4@���qڝ[x��:!�NaA���_�*���3j�g]���r�*�a{���I%1s� �\~GL��c2�)� @��-5ʻH`P�qd�� 낂���E�L��}��W		𿙳�c9�UA/B����3຀`������A�+Wn��DFF�^VUm�?��	��U%%�����i���^ 
1Ԧ[܍�ٞ��@� �Ԭ������g���:ǂw�Y1����6y� ��5����]#x�~��A	��K-���P��t]}��t_�Ns��ρ�|�JV�0�D�����@�O������6��M�J�DP7��'�B�k�Q����Q��H �_�Q1�@GVU�;�ׁD���:	'�\�G�(�^�O9�~��D<	j^�|đ[�����j#0���U����ٌ�P�!0������eho�eHp���y�j����~C�Z�q�� @s /�7�.s�'k�kHOK����~{5��X�g?	�`�4~�� ,�']�l��q!(m��~꺪��g���<�����ׯϜ?_t7Z���
z7�Cڸ���d4멯/s���d��4k��	�֣˷;8������<�Ĳ��g>vg�;�:��a���2�.�=����#�˗3;��E�/\�|���
'� ��w&�QVq۔�j����Z����S�tQ�N���׎��y�3h�@\���d���v4�˃�n�]�߆�?s��Z��g�(��*��?��ϐ���7�oKA� ��Ѿ���#8�0~|Sf7[���,�~o���w,m�QCY��(E��g�����FG`J[c��4v�1m�5+U)tN(��|��֋�ڛ��P�����ձ���*'��h�<�Y�G��/�ߔ)�(�G��Wb�{����3�j�Ӵ�YRt$�aЗ���T5�h�$[�^�}���7�f�TY�eo#8�h��%.�K�t�9ٴR�1��x����z���9�a/��GM��3�9�؊���+�8�V/?#)Q�9"�S���D"��X~�t}���q<�C%*������(�f:������MOOo����6��/�T��JKKn";�m�Z�����3�t���~�J4n\�X>�	�!7���p�r��$.�L��u�k ]�VwP=p�'
!�������H�:9>�w=U���G�l|�I;�oY�&�^;�����ˍ���� ^��i�v���7��`0�l�XT��!@XD�f�8�m�0�Mu�x�ML�@uZ���Z��C8�Șiܯ���3jB��TM���b�V��I;�,�ö����L��c��uc3Z��%@�C�TL�
�P�Ĥ��<ΐU6��ĹҰ�H��{͗�!���\��љ���S8��r怣�Y�P=$
��7{V;�9B������ t����C��s=��~��&z*�l�p	�#��'Xv����^���'6cS�9@�Lk3���9V����<$&�n7Z&>�}��.B�0��W":r.�1���F��"՘;�FˤLȳS���h'�NՖ����>ק~��:#7��8�Y�|�#��؏'��S�C��n�3u�AYV�C�&��v/�N L���뛙ͺ��PjÅ���W�&�@"�O~��j<�~��s�)#����!/<7�6�@}��-����� �M� ��Y]W�,d���nc�:C��@s #s5�����M�M0�	ҳg�Q�PW����ꍌXs�[�v��L����e�3�������"�`����ٿ�ĥ���|�^KSU�7N�Z���5((�)����?�0��moWF��'?b������%��$n�q+�z����C<P���e�õ�����}��F�~)��
$<5�ŋ�O�91�+�jA ��~�Ձ��"�l���\���:d���Zl`/�����/������޳����@�+����\��`1�_�̄�pc}5�AC��爙�m���6���i��/cx��is�j}��ky���)	!�a-x�$ԋ��k>�z��%j��ުS:4�pB%k�� "!!aiuei:~�&LEeOG�ZX0��� ���_��@�<yb���G����!��&b��awf���X���܊S��S�b��KR��)� T�x"���dTF� �>b{�M����֡ͽ$R�E�H�k�q];<
$�	��e�/i��X�=�kq�^Zs�����_�3�-f3���m^뺝l ;@�/���~���w��xrvD�sy�ZG�;�&&& ![�{]ʇ�К1�	+�~�fD̘���藪�$����\�)��?��Q��5(j�K�!�n�i�p-���ˁ��ƥ�S#]n�S�<~��͎�v��
��¸����s�b����9}r����_#o��YV��/�=� @��b�K1��4Ϩ����aI2�.�ʄL���~�.p��9nj`~.���_`Y�`���^�a.v��YX޺0td�)�1\7N�	�~�5����0eO+Ld7{i�z�+�;�4.��"�e\T�ub�o��������)�=�ů��E���`�����9����p�}��@�sy�'�=���;]$f���f�(��|��)��T�
�_��m�#�v<�ي���aX���O�P&T�,?M�g��.8�n`�?{D���cf?��.��y��Pw���_�S�-���U�C�<��M3��؁��o&�S��l�\�������|��� 
P&�R�@���`xv��9�L�^�j��4��kl���X��'��tEFs��]W�dv#�ƒ�E����C�q
�>$��������y��.�[���s/�zJ����w?|	i�ܶ�G=T�/�~/hQG@��ʂG�ϞH�l����?
� uCX�C@>�����H8����mm�w~X���Q�	��o���f,G�փ�����8ÁgS��뮀�Re��!wʤ*U���U�d�'�~����q���(�<���7����g�j�[�N����NX��
�}�����t���z�M�6nz�f�|��2�x<�!�EKϨ���]\�ݵ����j�5\d`/@���Æ���A7Qkk3fPq6�f�C}�ϡ��B�/C�G��:����H�����yj>�\�������
�f��C�,qf���P=N�^)?��@1SPy,k����i��CJ)��:]�	�}��%I�aLS�nZyU2�^c��k�/���}��������J�P���t�_�{���\mv�]���K�rgY����(��R��H{X|g��2�N�K@jXW���XI�	n,�n��������zf_>u^�}bN3�G����J�����20���O��l!����ƃt7ˊntww���xƐ3���{..2���V������^��W~i��1*�����?~\.c�ӌ����}<�8H�Edd����w:�1�}��ܾ��#�bﱟ��EB� n��%�bTC|��Ѣ�}nf"��]��+��8'������fև�K���U�pch$d^�UD�>q%i"���P�����}��pHto��C��\�/�鯫n�w�Z11��JTN�|�uc�#u��/.E>��ˢ�����a�!p4��#�4p8�e��l3�Ɍ',LOO{�S��ٗ�\�y�\f���]��x�Uz��+t�z����)1j��Цd2�\���i��v cπ�w�Y��"�J����
7�М.hλ����|���DϖP�����������#��� 0`�'+I�?����1?���nsQ�l�[�W3��y� ��߸q�l��#}�$(ˎqMʶm���R�������Y�mR�vp�ioN���}9����ǫW�~����p�8��ˡ�=\#�3����Ƈ����Kԓ����2ǉ��:ũ�N��}�xN�ߜ�V�l�q6��5��Ά�U���]$>8�����s��mLa6e������ 
�����)�۳g����c�aX�9٬pvv�3�)�mk㵩����{�Q&-���LK�g�ka�3 δ��R#��BT��T�o�b���4���@��-�_�1E�g����w-��;��9jZ�N�F��e>l�b�?�Vw���f}�9 ��=�Q��3ý���Y��+&^��F'7���|K��\	���Z>ˠ�*άn{�����CY�ǻk�|�o��2���R�_B����E`t���w������]�O� ���]�d��+�W�pZ�3�I���#d�������W�0� �^��ō
�z£3���b�������K��0�[��w���}�����W��:��7���8�5#�3�n���GO8e�X�ۍiǶ�P���#'N�H�ԖPn� =����0$����o���Ϝ��>�#���\%�"�<���T��׊	%�7�������T�UWo-**
_��� �1333�a����Qn2��GC����X)�;w�|��EԶ�<�^����ge�����b��<����<��ێ�'QWF�5뭌�̓�߄GEFU���V7t���1����a�UR�Qז��͎'���b?,$�d�8�hǈ' =~���[��5�J1�)?R��,@�+�"�UMS�ה:�Gj�O�x��|�n��x�i"�O��b����n2?�=,*�b�f�}�]0�3���f�r*�Ң�30��LO.�����������:�t��OF�=����8���s[�v�/8?_] ��ҙ�hl�<#Z]YɄŵ�
iii�x��� ����?�)f}Wz�D�^a�*2uNtn�b蛦�w�20E�DU�N����-x�Nî�����N�lV�b����啨S��qP$�r�gZ�������� ��/��il��n2:1��׊�>��[{"BA8���l<l�aVVV����[���Ш�����y����	�A�@1��Q�M�RF� ��J�6<_�zv5����	��E���~� ��@��P[�,(8	�U��	���Err��N��i��R0w������ˊmQ���|�ÿ��u���se��©ٍUY��MȔ\�j�,2q��z������O�C=��m'g;��K����]Ij��S<9]��Σs�*:�h��/��H]��N��v�P���ÍKH����R'����9�Jo�8a֫Py+����J�(^R?��g��Km���=D]��i�wK�����=��BMx�iݺuq��'�}�w,$��2>*{|�o�n*+��y!𾿿?��^3�>�t�F��N����t�q���K��oH��ܸ\�0@�Qg�?��E�盪[=҅{VX\�'��)[�I�[c����r����]�^?4T�l���-����>��L�Х��c��:��J�ˤ[Uo�z���w&�rܘ۾�i��ֲB��"JlL�������t��GT�z�.`!���x��I�m�9�wRn�ō��QWN�����L�޽y��A*����q�n��VT��C�\h��f�!b��'��!r�"mGݨ��7;��3�:ϯF��
��d�a,�$PĂ�{�F�7�O�RMt���渭�[F��y��VP~xf�	 ��{St�u.�ݼy���z��v<)p��QZnE�7� ����A;�����eJ�=z0%���8�����������cc=���9�Y~��]��@�����{w��IWq�ؖ���y����H>�	��	���ު(̊W����Xu�u��?oK�@�Jʚ�9 �w0���W��ek(�}㼼�Zx�3�s�n���_ܷ��w����ϟ�X�K�������U�`a�S{H&�''|�_I<|H=K��իxH�E	���Snge�%��g�]���R�;���K�Q˴N=z&*l��w����׵��B����f;5�O�x^0��]ӫ����oRX~lY
���p��Q��'Oᰜ�@~c���G�wv ��9k�D��@�>	�K#<4�A�C@���-<��q(R֎�#NM����2J�����fx�4�-�Hr�����S.��T3Ѯ�y���K�>�zeB�&�g"��0�	lO�=z��)MM̓J��$������^�O��o����2aݺ�1��?[��Uu����C�%P���p�����G�3�B1e�?0�a^^� 0����o=�J�Zu��ƻ��H=Dp[խ1�6���\\����}i��J�g~܃?�p���s�#�2g=Z���� ,�q��@����BɒkVPٽ�!�J%z�K����ȴ�
{/wR飝���?����w����]��*W����U���w����]��V�8_�V�����A����׎$�OLW����ΩǤ��4�+�61P��������$�_j��K_��@�ܕ��-ZMG������w��+�]���
y���!\����+�]��
W�������w��?Vh���@zL_����=a��pqպ�߈"��M�-��IwB~�����G�p�o]߉�)}���1i��� PK   ���X+���  D�  /   images/5cebb09a-e86f-4cb2-800e-22da09d26481.png�yTSW7k+u Z�	�5�����dK+�т*�"�2$�!L�
���QF��bŀ"�@ ��IH��D÷Ͻqx�����w��ֳl�9g����>7湴��Dz��EA���k�6�������o��*���>?���=�'|^H�{؇@��A��W{j�<\s�W۳6d׳�c�.*��v������E���/�_K l �~�i�����n?=~�d��y�>����g{�.߱�k?����n��������k=.����yAʶ�S?7/ot�Qi�y�u�̿�]1�����_y�͜�~��z;f��ln��	�	��To��*���w�y{YJ��|���\�wr�k�0�g��2)��@�0��P7`2E��]��Su����\�64��b�BU�c�C�qs7E
{�U����|�
d� d��\�դ<M>��ᖼ# ,��m���/;K�5������k*�pnyv����ßM�GV�m�o����߆�6����m��m�����	�(e֚�ܩ�wW�^d�����RX6�,H$}� �o�h��x���X��p͎�Q���cNKCnBI�q�=qHi�e�{O�1=
x�k��U���m�n�$[G��3(��S����(WX�}�O��	��@p�9r_�6���9m|!�X!?��5>B?k��9���<W{���z��˿`��o�_� �ix�2������{�7��k��{����W��r����BE�z���V���7/��e:�I�ېc��2�?�)N�oL	G

�������/�O����"���<�Ot�"�<��,�z瓂]ǿ�ϡ.K��l�V)�8K>/��i|bH�	��w���*���w\ &�[��F��Ld��4�2��f@O���Ӛ�h^�d�+��K�������	(��S�|M��;) ������F�gAB2/	?��{��8y��v�BX�-���"]CY�����i{�\���D�=��j0���f�/q��!������M�u��>��)I�d��dK�nɁ_����Xދ�9s-0`�R�c8�@@�5����5�/$P�]�ر� �tZ�J�+R*9��|@\��5��v?��>���:��:���$2����Lb�z\G9��~\��.'�ny��!��-�q1Ș|B���_]$���	������|oS X&p�mW�c��~�?���{@�9�(���uX�MH�-�0P
����`����$/�������1��1F ����7r)D�v�s��Z|;�\h�D,1W8���gƚ���8f|��J���W���~!Řn�ŵu<��K|���ޔN�]�.�v-��r��7mrue�'q��L)R��+��¥�����z��ϑ�g҄DM�f*�r�Trܒ"S�+�#�+����ϝ��f!(7@?���9�#�?�}�+�a��כ�+��EL��\��&�I��}����I��]��g\B��Xe������)=PI�Bc��<�p��Kb�DB|~_��[$� �Q��=��g�����I2�uC����,�=0�����霫�3h�����tG��n��!�Y�^�&��~��"}d�}vxf�=<���:�G� 1��3���`�}n�ϴu+/?_��nF�޵��D��x9��k��K�n�i��+�0qa��1�y�8��h5Wb�م$59��C4����.��9��ӀT'ɛ�<�T�/�'6����~�򼚄��)�YT�\�	���)���/(�Ye�� ~��J]��*����-M��3H1�nlش-�{	0�`{7i�$�d陼'��K��R����ԣ�����]�QG��P.N���2��;��/��~%�mRN?f��
���<�WE�s-t 
��v�Q�`��m���4@FfUyrv?�m�))������-�����2.nxJ�Ǟ��߀^OJ���X4F�M 
�m%	maz��k�j���O��� l��fI_6.;�G)E=ΫM���/N���쳰,F�Z �z؅�n��?؁��< ��S���¤�h��Ge l4������,�nY)����i���8���>c�7����x&|Ό~LNߖU\��*��9.�S��(�5����^����@�Wǯ�*�Pq��R��ySL
����oâ�z�T@�� �ǯk�.�)�kD�G�e4o�����o���UT%+?5�DO�/�pƁ4����}��"�sS�b,�B5�/X�ٛ@Gr��!y�6��ē�M8�7�I U��� ��[Z��B+j��t�|�2s��R��I����;v���Eʢ:d��ЙT��ob���l�}/!�0�_P�u�[��gߊ2Fu�܂Y��.�T�����f�>�g�?�nY�������g��Q���D��R}=ax(�^~��?06����G/�v����p}�37���o�����s�"e��X�����z�l��cZ/�)<�u,D�Sܮ�E$ �CWL��U{��� DC/@���PcA3��$Z��{7�(����a�]*'��� ��̛FP	�g�G��S]D#=�
}V��.=�칵oL�\gɤ��Ìl2ܚ��N���i��6@KI��7U�>W��ʷ=�i]����Y�ݓM��[�{���ީ˕�ח�>H�=/@��kg��4�|*πTYU/n2
9��֕��^H����.̥OL��&�I���{����]��Ш��k�y[���X���d*���D؆-.*��}�l�U� ���Q����l�e��e,?��b]D~^60V��4���Ӏa�̟�SB���py1�OT�78���-ߎ�5����Dx~ء�,>@�jeSҼ���������rt*�s�!�[ͧΊ/S�F��x2�A�G9P�GT�� ˞��@���'��F�L�W1�u�p�X��YAR[,��8'�$ 2����0��o�=�
		Z�/�dvWC�O���{���.Y�4w<Yw� �Ke[�v����˝���Y�Lw��^��5oW[����e� 5����a���r�/��Rq/��.!�kV�����#��W7�h����S��k�|�Ю���)V����<+KbP��i�,2t�=7�����,g�r�S�4�՝j؝�&���X{L��^�͝�H�����浺K��,=t����O=��`=�k�i3A��xM�t�y��W��^�����O�gﱦ&��~M�pG�3a��f@3H��qo�[΁���ﾡOm%�Z���53�9o�,E�aXĿ/����Bx�_f��;>�B6����M-'�x(���];��k6*3�y��"�ץպ^��r��r8e:��M��%��G�F��E�Yӯ&گ����/�Uk�_祻����}I��hi���2o��6�^��_7U0���p�<��%�?LD����л����g(������ ~O�./o?r�}��y�3��Z:V	B6��U��3A�u��ʨd�jD���\�Κ����ӓGv��n$�[�l�} Ȉ��H�H�m�O[ó�3MI�n�Y~X�������F�A�	5�h*���U�k*�B+�7�Ŕ�(����YY�ɩL8d*Æ9ߦ}Z0A�O���N�'���r���Y9S��wnC+q�������2�>��N��R�5y{!wK��(��x�Ӏut6�^�d�_&őo;S�M�wQ���}傘ۗ�v��?�����=�2�ϛ�J2A<�#��nV�x�[��� ���]�9�]��z���,�:���Llʖ;��� T��3&�_����^T����2ET��q��N����9}�O$�[��v� �͕�,Q�̶?��܂�Qp.��8��uE�B�%5�X��nb�W��j���MY�"���U?~ j'�rA����p��&�7��,�0�Χ�K�P��sE~�*�ơ��r����ͬ�?�Q�i7��̏��:8�H�2�9/l�(H<����^��#�$;�G�z\���,��t��իޗTV5���^���l���|ϝ1����v3�[�9+�je�ŕAc��hk��R�����'@�h���FM��m�	[�b��`��baW�a=�((��2�or'�T�9�pZ����]X��,+.ˍs@+�{e
V�K�n�J�5(�0��P�$K�Գ4z�����wK��nO,!,�N����k��SE�j_��ƞ����z20�kT�l�3������}�{���R�A/=&n�b}�k���8����f��YŎ��DU�?��n�����䐻~ؘR� �j�[e4�;:�ye$"�C�w(R�3�o��9���{���=��:�6"��x��
k3������Ṗ�ɑ#p���ͫ���?12�^m���'t��2A�f1��Rf�M��h�	�D�:[�����h�:���p��>E�JuY�p�*Cʇ��;�`JLz�4�e:2������˗Fb<�f��+��J�W�UG%'����j�����Âq�l�_�τt��@ς4�A�5��|߄�v����61��Ϲ+7�[�,���Ώ.�����}5XA�)�X���ޖ��4TMWу��d�2?3.� j�!�9���~+n���rM�MG�#Z$/�¢	cd��6�}�d	��ȟSd:1��l3fN� �d*O�B�f�sC��g��<�}�=�����^��Ct���]�'��$d'�IcZ�3�ӧ鑓��nر��؊@*��i�5YyrJ.]�2$��1?��WJ6��C�xoz�qxO��-^�˭^>���U��d2�!��ݿ��5�i�իF�'��:�fBWE�撈����s#6s��:!�Xh���R�!4o����I�g��5���޾oW��"�����(>��F��=,O&��
�ݱ9��4(�t6���8��kO��}��l�뚖���B�T�@�I�|�>}d*�HUd9*�9�p�ԂE����7�^>�z�u��m7�7��;8��ksD��%����B�Cy�90�0ϲd<ռ�X��A�3�v>{��1�aEw$=�%&�S�o�:mW�b�:zs�LNc��j+����c��e��O@H�Xi�8��c� �W�$g�9�#����1÷o��&r�A�.��j��=g��MV�tSjy����ѼC�F�/�b�Q�W�@��Gy�"�Vrzώ��Y���*�6]#V�a�G���nP�^熯fl�(ǻ %��!`K�����"�{jd�Zw�8��xr�����
,����?�ԓho�F�rwc�4�c��Lb+��F�P0�[��2�P������M�����>z��|�N)OJ�eM����7�E!v�6�S�̕�#�;�/�q��쌺��}��Y�v,p�W�d�R��F��x�_�V8+Qm�WD��>X�*�wI��R��\ϭ�}𺎌c�Mu��2��c���n�L�;�������HQ�Ik�mS������ғ��*O������:���d�oE� �OǷ��'?�gd2��[�^���3�*i��lk�G���F�҃S�\�G�L��&�ۻ��u) v��h��f��+�T�����o�"F�_�ʤO�	AP�v����<�9:�wk���K�=�X���@�ުN��{��`X+JP5���ϳ���F�9?�U��a�4�R��m���f2P��Aek�0]�"z?�8��044����t��s���93�}��'bz��!NB��[e�zN���X��7"߂NaY�I*�Vj�c��i38������0�ct*���4��s�J��a�ݮsq��'��}�3���vO����C�BJH�LIP1�*OO��ARt�oc�յg&��X�EO��}����%C��dD�Xi�ዪI�|�lK�ڷg�sĺW�1���S,�xk ,X���,c�ޥŦ�c��K��=����a�}���4Y�v���T��2>��7�KX�iD�
NV��ED��02S#u=�*���Ao5���� :9�/t�����u������}K/��5��y���U�L�mt�>�K�5��'ℸ�N4'3uYc�d�г��H�rAv����9G�0�
y6�he���:��l�Z���?l�\��1�R�a'õ�(�������-WD8��̅�8p�s����dQ��-���G(����5o�����Qf��]n�"��p�7q��:g�H���?YK4i���]�4dQ�ץ��U1<��;�G@�d�x�_�6_M���'�V���r�e�����_���#_,�i���5�N��YGWR��?�O�ׁIVeW�9F�s�<mo�#\���&e��p�W�^���ź8�5��כ���CR+$���k��y��nWx�p��S�i�����7n���A�g�X�{���g��5j�����C��	")x���H$���[+%됐M����i]�%�q�j�>iꭠsނ�<��HV��OY�f�#$d,H�} On���Y��� ;g����U�ae�,�A�"�I��՝���"��ꉋD^�6�;�_zeF*��r� ���P�9�{��� L�F�$�h	�G�N/VH������%��I�^A� ь3>%9���^�;��&D(O^Ȓ�����x�,%iis�������?�elb�5Z`�]]u�[�k�N4�YwR�I�k6�Yp�C�%����$"i�u�����G��?��ҷ[lւW|���. ����Y)G�6�w�/��>�b��5�1�k��IY�#�svA3��~3��5�'�3@�_�e��!�G����iI/�d�O�
�w���j5�	�~�����'B��:�g�gB�;�u+��+Wʽ����T��%����ol�q{!~n�E=Jv���(��۽tٗk�:Bo�^�~o�*"�mL�W ���l������z�0_��ܻC�̛!z�sn��iV�C$3�Q��!f�+ -�ˁ[�d�Y���|�FS����7�����Ր�>��vv[(�l��A)ØL*�]�������&��xRnC�"]N8�N#F/�;���d�,x�B��M��Mi����M5w���(�p����ղnR�뒧U�+yD���::|,Zv.�h�ic6ȱ��v/�(��z]7�����F�F�}N�U����A=ą�Xaӝ�J6������=d\�����-��W���x�]�A.�-�1��p��Fr��-n�0Hb�Ͻ���e=��XԀ�|+&+ł{84�<�6�Q>�#`�m�3g��l���G!�Q�U?�e]o��{���@��a�+�e�p�)	�L��ҋb�1c���0�<�'���=�I��뾥����;����^��U�ǖ@��U��О�,'q���k��t�J� � 6���r�v��6 �O�&�+lm� �lTvqb.�s���|�<�����"+�Y'���>�W\�o@��0Cu�[�d1����<������q0b�����-��?��Ϗ�E���
�W_���ui��(܅��"��]�n��
��Ћ(&�/5U}� ���?��Z�?��̙.jP7J�}3�x�ţ�طKlA��m6�9ѼK��d+��6l:k/��hE67ѝ�����QY+��6ő�_��MK��_e�_��Q���j,����+i��<"@>���P��R�t?<wφ��L|UkV�	Q�Fу$^# w沼]���CJ]�Qy�U�U�	�Tͱ�>f�=���J_���~�e�m����Q(��Л��å*#d�)�e��8q�7��[lϕV����b\���%�s �"���/�:L���B�ܣǏߓ��:xj��>��_�?���Ri2�W�&�|�֖<\H)0FGy*#p;�xq��TE?fj��$"�����#
L��|�et��4�
E�zص�f���;k�ʦ��yy@�a�����"��X��y6���	�,:9������̼��h^|83C*���'
Qc�˝ԃ<�S��W�Tp�d89JL���#sޯ�C��Y�G�_���C�Å{'���!g���Wa>PӒ[!7�Τk[�s��	Ǆ31ѣ�%� r�4"֖�%P}3�4wo�@!OzSn�t�?jۦ"��!`�U;�Hٺ,�r3'���y��6���k*�Ȑ����� �N�����o��*?��V�K����&���"2�>=2������x�ꂝ�:�'����T:Q���{�i�s���;!*�ź���2;;a�E�>8���tV(y���S�#�v�N-�Z�:�7O� ���E��I,�ԆUN>5��n�U�١��F�w�����s��Q�����'|�r��l 9\�=�]y�5�c=�YsK$�N��0��݋���ħkn���B"y�77W��ߘF��2
�,i�5ֆ�*���Z�*�<߄��0}�Rcc<=S��M_�c�y��U$�e��v�}�����4,�ϻ�ɒ�pB��c�u��+ƶcw�̀]oKQ��ȱOUQ��d�Б�/�5O�N��O�.V��ѯ���簯28�Ra�Lb��ֽ���W�d�*#2��+{�+h��u��g�!y#��;����h�#�Q̖4<׌
F.z-we�>�]D�)j[,2a�0S,�����"�8��������)t�;����8�	�J�ؤ'�{���84��{��4�X�:u}����@�7�`U�2[�7F/��/��,|�M缀�F"uK���x�Q���� @0�Ǭ���2K9��Tj*���V�{R�!�X���Y��{Fr�}������҂9��z����*m��'V�u&O���07C��`n3|Q�JOQI��L%�᧥t�~�H*`��Ah��~'�߃`0���Eu�Ƨ1��v��B�y�l� ���v������Ij��&���:��V �AV�D�P�Kb�2��z�"9$�����#�l����T����EZt��n�:�O�0h�W���\}!�W��*�mXA��@r�0������߻���,B߳��G��P��\�U��_���ܝQ�p���Q(�LuF�1];��'��WEK��M�u��� �o�Zՠ`��=tt�&-�o��w�k�b>��ԜPQ"�V��N����gY{��֧ؔ
ȧ�ﭜ��%�y�5�LNe޻Lbx�M����V��qs�������Ѯ�۫,�Xюcok�$/�����'s��3T�R��Nx��Z��<2w��һe4��G�᨜����JWE�z&o���ס������<u�-g~�S�w�D	�����'	(�Mb�2np8�x�v��@|fO��NM8�'�9�Ei����u�f�\u.���u����M�c0L��3���\�\��aw*��~&5�`��`&�X}Q�@��)�ܰ=�J�m�b/�-?�f$Ɇ�є�SYVg��5�V�Ƨ����	�����T��W���ط��9�^K��\����7q�L��TqWS�0�9��]��6��~f���/���t�"":��.I"�dl�[�J$��pd����q�b;��[O���&Z<׭���&���\�L<�\�>@ՓG��O�mﮬ,��7���Ń�r��L�mFb�X��n�+�L}:�e5��7]�]k��u��;��������78��M��A��(�~0������M\��׎WaZ��?�k�C����%�S�������j�\� �e.�A�ͷ�KN�^_�?�0�l,ۊ���?4l��;��s�������c�!ǖ>������W���46�d%%���6F�M�?�=�&��GJ��{�%���m� oY�+u��%�2���ލB���O��1/�,B~�8>V�ܡ�kVZ����y�I�jnk����!�Wu���Ti�l��nz��Z��UUAe|���T�iw1�����ޞ�&��G���@�W0OltUb^Pc�0�;̺���:#kC���ix�f@��&�um��1H��������$� `�&'CrP����	����4QPn��14;�1�<��w�;'�e�=�`��y-�����-�o7#� �\�r�i��b�� I��b����eD�W5��;9�s�����EF�GM�� ����#� �苩F���w�\%�����.�5	y-����l��i�B�(�YQ�� ;�c�����l�bu�ȿݾ��Ǯ���t׼W�s[o�m�J
���G�6��Z*���EZ�BάS�%%	N("�}gN���iCEW����J�O�c6��iK ��E-�����|�P?�H�%�$_ѺoH�w!w_�R5�!s�'��M�:�&��`�D���VG8�$��{ �'����B���W�.m��x��&�T�3�I��)�ÊHg�;>X��/�M�
��7���Wj�[����AE���`}�${���DG �����]��j,E"�����}:�R��ԡM8��w;X#������]�g�Jb%�:dٺ	E��� �V�e-������M����z�����WM"zl0�$����V(�~��!S-f"e]�q��Asl �}R'łO08ZJ1ʣ
���^�h�����!�*���#�s�-��R�o�껡O��1��BS`��i�Z7\W�,�h�(z;Y�/(B�V����D����~��O��^�C����Jt��H��`��^�UZ�����A�vrHE��:��*�Zl��=F��] ��r97
�{(��80�U����׬���2+UQ�,(�dGlpn��Q�^k��V����7�)���B��Ƭ}��0�I��L_qBṄӃ0�!]���Q��<��)c4J�\D�ښY��
�]��{��&P~vR?�u�hf�/gw�>��6��e��i,y����O$�����?�6��Hx���7�۵�ՇYf�(;�Ʊkrb	��3І=��Ё���
�1�f�s�N�+y9nͬ=��jTTEh9gNs�:��Y�>��n /�rQ�`��ͺ�86Q�m�O��F(��,�abS֑��W����Z�2;�@�M��B�oL��WP�s���HkH��Ԙ/��]�;�)F��DA��w���ς4�R����>J���8I%vU�\��tY^���������T6=:@�貊<��ޤoD
�Q梲����=��\������Xw�n��yb��{��[S��X	��<Z.�-Uk
��h!�4Zχ3y�Fo��q�㎠G�[3�#���+m����r��g���5)��eu[���׍�O�{��˄��ǭk�H$N����=�h���SA�p���x,,���'�;�S��o�mIɕ8� ����^��I"*�
~�#��`�7�K(���Y�*AD���sީ:����B�Z0�K����~w�~w�� Ф2��{g;N���i>�g`Mm��d�~�������W�޹K��2n�Qb3<����687��v!�Ȋ�nǤ��(����@�W`ʸ6���ŕjl3��U�����W���q�*(+z�C���^�I)1��iQ�,��9S�����7����?�6�iJ�L&���l.���J ��IjB]��Õ��,�0q�4�ĭ�3�.-��������ae
DX���$�-ޔ����^��&���Bsu?�Wʦ˂�a�ll��Z��vL�i����}��J|,���?,;UA��DW���^%E/���/ l [Z(��h~d�=7��1�zN;%���u^KR����>�;d&�S�UVi-���xlJBW��S.�1��NUR�s��9�'Z�C�F���$��O��M�$��V!�jeEH��9��VHܲ�%E���[2�nR�ʈ�w��	@4b�����a�>�n�hY1�$y[�>�����V��$�!�$QBv�2�2A�rkT	�!	��Zx�v��W��W�f٤{O��l�,��������M{�X��z��T=������f,�}��Vc�/]Tb���	"��O6.���nv�4v�93��m�H����O;�7(MBR�u��?2҆+�w9��`���x��T����z���n�bk��m���}����v��`�}km�+�HP��ڵ��mbW,�ųQK����VΤdطC�~�1�й�z�u��2��#u|p��c�E
�L�9@磝_m��!2씵�s�7ǒŋWA���n�qw#��,x?����t�N�}�TF�pi������A��U��ʳ�74s��g��o�	R�D��R��]+
�3�}v�vG�.�KRTl���D�:77{��)�w�<~��j]Z.Ҋݚ0�t���^�^�"zd����	�������k��F0UdY1Ɇ~�>���p�|�b���R�goRv�R��R�h^$˗2��6�ȳ��RQ�س2�L�0�_��l�*��|tW��E#�S�ÞX�:����#�!ǆF��Vwl��&��[��uqd�x��kU�Rk�m��1�W`�ˊ��eww�E${`&隧/��	+zm��${Qa��A��qTζ�߿��Д9��*9����'gH�_��@���>����"Tb��E �U��܇�J������#M���D�3f�3$�y):�O�qh"F�lo�5�(�� �{wD�PK;q��7fN�@{���h��첏ަx�TO�&�So�;��_�����[�L&aP_ҰP$���{��p�E�fr<Eg�x�VT���]l��D�����V�z4;��pi�bѲO������dβ^�w��{�hrm�(e˧^�ٻ�r���B�7S�~Is�I�fό����{oH�ʵ0[���?4(y Z�b~��m].ت*�"|�����C74]��Sf�ZB��Ѡ��j���w�7Hϑ�`	���=�7���e�
*-�H�l�l�P��}|��|��ݽ�c4w���]�e�e��3V	�S�d��������������U�gz�w�o����S�ߕ�C"��?m_~�F(3FlF�9��{��Bf#��� 7�_D]]�km�/N� ��G�����5Kn$�M??X��,m�h���ǆ�#LQ�T"��$2u%��W��E�¼3;��%���O�>�}�]��Q��k��rU�w�~�ݿԠ#�Cm�&�΀�gb�B�N�ޤ;�����
����+9��)�T]:��pt?	E�q؈?]l؋?�!��y�/ߛ0TT�c/���^9
�����R�5�n�ry1Mcǩr�z~,>��u�(7@���.���>>�.�>dﻁ�s�A��ό������;GN7�I���x���(����f�0|�Z����6��tP�d+�9��޼��`1"���_t�[���	N��-�a�ￗ�?*��i!At7< �_���C��"#����6�(��Ձa�o��,K�#�b�_� �s�P���&^ V���� J�R�8�?.��n_�D�
D���h[����{�W���[���h�J�*��Կ��9x��P>��-\��rMΨg�,�~�g�$^YG�@���4d�(�g:�@��O2���8S� ߳���ë��9]�L�=��C�Ps�>%#���w�h�VV�$��p���ҏ���ύ�����[:E�g�A��qf�f���}���ݧB��� b�@t��;2�b����m�'���e��Vf����C/e�S<���B�p��`����'�ϋT]����i�y���+J��X=�:1�������6LG�?+��ڗ7���p�QL=�|�-�6~�Sa�}����?h��qh,[���T�S�QW���Pg��|~�'�ʣ�J�������q�M�I�c����L/�]y��������ǣ�K�ZxIk���'/�����'�g������ߔX_��&Z�Mkwu�i9�;s�JMG�K��3�{}&�EcZ�˃��	󗲏��v=Z?X3���x�7�o	B~����d����fvK�o�*���n[��R����29�4����df6�hl���r�14����	����'�(�L�sm��:�&�l��it������k����v�W.�|�,1:@�y󻚊�[hY/ð:}�k�m�ua�r�ע�\Ӽ�O,]xb>KM�͸ߘ>�qg��4��aW�;S��nq����ܾ��6��D�H�Tu��F�*�_��sA|��N�o�.��.�!!��;��LrI��� ���q�B��ɺ ���<u�D��<ǘ����"_
~`�>�'"H˭c�e�$G�W�0)�Ȭ�������<Öz�u�����Cu3мΰ1�Ÿn��5���笍���Ź�h���w�\s<�v��C���_(�]1!3�U����nv���=~�����b,EU�
�cDg�
cIP��"���<�Z�Yu����½JN*7���|�$�Pr��1N�����\, ���^������4X�ZO[k\7~����cT��|��{n"4�v�I�'�'�����ĉpn0e��y���XP����x>��Q���qi�/Ђ����d�Uv��k!�_I�kj�?���)xH7_¹S\ëU��`��\�p����#/�Eg��n1X��3�e�ck��ԉ��f�gic6��.ٟ2݉�����]����7�(k+���S�l�fΐ��f���s�N����	gh.�c��޸h/�B��v�s��WBw|ǾU���Sx�h,%j�^��~g��Ժ�`ڃaRlͅ2��;D}p��������ɡ���>��.�,F�v�)�K�i�b�%|��Q�2e�f��	�z���1�������r�DO�@��.Ɲ�Q�/����⿭	��}x��nni���lY�*N�	����]4�pt.e��3�/!���(V/��n:�R��X����1�K�����#����B,G��d�`MP����4CO�E��C�
����J�6D��&�{7�������pc���4v�(%���+�Ldx
��^	f��,V&�^�{ɸ����ע+'8.�f�ܤ;K �~�Wf�}�W�g/4�;KQ���[�RH� o����<�>��c��H���u����o�d߳C������N]A�P3#�D���'�A찌�������W����]����Pa=_hh4nf���I�`�Zh�ë�+������nC�>+�н�?U��C���N"c��JpZ�5u0�Ĉ�(�1���+�*Wxx�g�׽�A�Y�Ln���K��K�N�i����`��^rd,V��[%��ĕ	�串>��p���)8>5��~-��`�[��_(R!�!Y�G�j��.�
�������&lдzq�P�������H&�zЕ�l*��o�V���B�W��@����W? i�D�ME�A���*���9����T��U���u�ش<�B�	��'��hT���tV��%m�0w� U�� n�	�²��:lΰ6��}�>��Jc��P-�趁ƓPQ��j��24;<�쿁����Y�uN� �6�n2L|��c�Ze�������OyJ�I���u"�c�N�aϸ��W���
�,�(�Qe��9�_=�7�����X�	9��������r��w��o���R����)�ܥ@x�z���J̐uxn���>�&�«��_���Q���)�T_'�����,d��sDK>����zv�ܛ�n��s�!ӱ���V�Pgr�����b���\1u���*������E)�A������ȹ�öZ�v�
�wc~�����x�jpY����G��]Y��5ٓ���=�dӒ��#A�_�gWʻ����p�\�=�~��[�B��xZ_#��\;�局T� 𭀓�mr����;��"w3Ȇ�&����G�{�Κ��vS6�=��!�D4�uY��8ס�/8
�Bk�ˀ�"i�C�e}��M1z73A|Mf��ҰY�z�@y��nc��~�¶� �ڟe�o��<s�|Cs*����r���"�۷^tS����3����&
��P�p��DHA�yj�'��W�َ�/��
R#S�F�t��b�MP�L�Ȭ����?�ݑM�%�>��B�-�����~�:��Y��CFݺ�'�FH��m/���&]�cK w�4L�������c ��:��� ����ox��� �c�l!#�}��χ{�<5YPk���
�&tU�������.*�O��*���0�����G2M��IPd���H��@g
�BJ�'V������d.��o$��=�V�H�{��9��--~���5��p�s<��OA��	�%=7�T����T�Q�v}v̄`"����i����.z�����UiJ�w��(«���q��� �a��]�*#+�Q-��Q���uZ��� m{�ؐ߉qة�i�������:(�*x�j�b�|&��;�_b �����豙9�R�����qx�a;a�추}����s=�{����x���4>��&�G�I����(t���v��$���?�J<A{춤�7��7��YH{��.HQ��y���O��_��قt�������6��%D���1��'E�	���]�
S���܃߹��?�Ci>4W�Cw���rg^��xڣ�v3P�*��LD3����������{>S�Z�ڙnX]��xb��s��Q�V�R	���a)�-�[y\����B��뒔�^��i�ِ=H��PX�
֣���/�|y�L0��#�h�ɁkWf��<�Fח(��SRj%�|�yø6��w���hc��=7����Z�Z��/���.|����Ԃp�-mݝ���:0=I (��D���5�Ѝ���#�Z&~x��_��)��`p`��&(Niݧ����w4��ܲ�o=��9�����TBͧ��o��_�� �Ss>�Z)&�+�Q��f@��VN|��i�a�D���w�A�~*�-%���f�q��] �㷂�uSw��2�ED�+���Rv4#���y�VD����s �`wu��Ai��ϱ�x�8^Tkx�B��&�=rө6Y�hH�P�F�YG�U�$�Z)����ۍ�.��gO����.��ʼϠ�5�7�͖2R�����k����n����?���T��=��h[]@�ր<68<5�y0���H}�a�ƿ6ȱf�����z���_����y�\c� ��:(�2r���/$�Vx0#���Y��ꚴȹ��� �:��q��\%,�|*%��.�_�S"5�����1�K�f����� ab�z�U�w|*�� �G8�u>+�?G�]�Х6H�)��/$H��hOp��tZT��Xj��Q�OQ�rȭ����z�~ss�|E&YF�m��}�R@)�3`�+��F��C���@�A���x�J������o��؉q��5��U�.A�,���O�8�����kL����u��tR�f�C�9�K����Y5Q��f��L�kf��%��,HF���'j?��(�+����JI{�����A^̪�:����>��'�E���Բ�SÉK�s������0���H�6ۏ7�/����=�~W*{�>�B�;z*�?5��zq�v���$UR����BZ�d*�S�(�E;���=�OL�`^�ߧ'%��A|[�V��‶��O�/��������>>h|�s�]3w�i�o�\9:m�&y*g�TПL��ܠа�4�M�v��&��lt�;��XP��f�a�j������t���X�r|$_�XR�3��y�A	~�k��I�˚��g�g0}���ᆪ>�ϝf��#��h���1�4�[9��.�,���c.q=�cQiD�"�:pݹ�Sr��u�6�3���n pD��DE��8)6rt����'�p5N���ظWt��ҹw�?A�6��ā=-�#��V[�>1Y��q�󠎼�Â����B�u����v�-�3��
I�r�Ӯ��[��*��F��#���@�~�x�P��R�/T�d�����10�=?�� �R�ٓ����I96.-271qH�.�vJ`·v&?��{�s2�����ʘ;XW��JR
���L�Qv1�>~8�B��\�9Z�38�Q 662��6����(.�c�\�|wV��y-��1n��8���G�e*��}b E�u}�������eϞ(�L�Cς�&�!��V�Д�tg�n���lĳ���,�EJ�YJ��v��J.���v�ƒzD�����P�q��<�w�|I$28gBf�o m�[���פ]f�P��l��ar�n�ׯ��-���ySnG������M�y5Z�xGZ]-�dP
<s��a��B������tZ�ݙ�w��x;�G��T;�R�`�dW�˧�ܮU�O�8T��i6���ߕ�)R���E��(ʺ�&�>����o�
��A̭�X%� �uϩ�<�)�Y���a��U��L
��a�:l7Q��Ɂ�y0���T�n�0E�����\����t#������k܏7��k'��K�j.ж����?�Q��E,�B}H����&���� 7!�C���ă���]��Etg���7;�)d�ڠ�"�K~I����E	���.C�l��,��@���;�����&����K�8�]Μ39�� ���~T��?��mOj*��hYMڴ��Z����(5���ff�i���7�߱���F���e�ܷ�;>1�����\5c+�_���l��eh�4-^�O�#��R;��MM��,��8_�HߺN���!`���8j��T��N�$��� ���WAk�Y�5�H4�M�u��Ű���������Kdlԁ��R���|-i��p	����4�x�q���O+��s��Ccq�،z8��T��h��3FpP��l-Rk`bbҎ_�VϢ9���~�ف*j�h]@��i�M�����j}3i��.�L�⍸ۆʒ��g���?R����
5�F��SŴS��G��&s�%�؍��[=jHڅׂ�f�%��`��:�V�(V�"8T�s�MA#l"�X谵f�hE�W�q��*`P3Y�:vtkr����x���RvxL��������Me[�����+�s�+2
�� ""J1b(�0#�:��A��Z0�6�U�Q�9�HW1 "E�^"�`��[B@HI�PB�w�s�}�?��|���|��>k���w���0�E ��b�>���f�}�J׌Ω혢H�����"�(�=;)�B�OG��h���[�ƾLÕ�[�i�e�6��!Ơ��LX'R�����L��*���#[ ���(i�@�M�Ǔ�lI����w����*It�2���_,�_qi�������w��_˪�峁˼(�+G|4G���>�5ޠ�Z�k�뎩��ʾA�6�IO��K� ���i�چh�S#1IJG��$�3����x��;�3�f�~�;�H��o�鿁3Lr����a;'�Ľ��X/tLU�:����N���+��A<����N��j�Hc"?jo��\[d	��mp��F12<0�67q"�b�%�)y���|�&���
l�ܨ=�լAY�B��M���M�Lg�OR�tZBC�5�W_��~B<�;�ݝ���oz�����z����K��i�m`��k��ȇhّ����� �a^h§��U��g��g{����7��������vz�ޚ'|��� a"�g���`����SV�L4�Z�b;��]�m�c	(T��г��l&L͛Z��V��݃ڪ��Y���zk}��+-��L�Qj�`��Us�����=4i*�ܴk�L�U�;��HC�Q�x�4Ӹ�O�<��w��ʑ%hr���HΛM̮�>% �䛚����Ԫ��	k�k#�3Ea���O��{q�~;�Q�0�-�J/V#{u�����K�}:�+�%vh���L_e����f���;n�(�3�f�F��W�����������Zx�BWؕ���f�of�q���Ӓ�I�v/n��[%՜/�ܨU4x���R���2�gO�.�G�R�p�ގ�q��)�6 �kY����$٣��#�/b˴_�k���c�������_����HTF��F�<cN�i	��e��� &r1�Cqdۼ�5n���J���7��ՠv�k]+4�_�q�ablxX"��Z�Y�m��uL�&1y��^�r<��Uk<NtZX@��e7������ͨ`�V'����˦ui'�xy}c�s.D�#.�@��U/�g��h�$c+ҋH wt;�2�n��U6� ����|���z���楳"i���3_U�a��ZV��\�Ò��K� ����v7jxdg����L��5�@�F��U�p/Y����ƍ�S�x�4���y�7�1�}�;�7�c�t��o�ε&Id��vSb����;�ƀy����x����ܐ��dgb�a����2Ȋ�[3%��W�v*�x��-�(����o'oC�ܷf��M��N���!�ԥ�YX��")��f�w�:�e���r�pc5�#�a��������u��8R^0lQ��ޮ����>8)H5T)G7m�
5�o����3y�aQk3c���#��&�gw5*�3a��S�޾���Uʈ�a��S6;�[��ns�@U�Bgc�����EbXf�� ���jO��[|%ju{Be�W >P��p�V�G�[;/s����*)]o�>������aL[y�
����{���4�s$AK����c���g*���Ab����TI3�$���$v���.���x�Ǉq����j�"�X�&;�Z���1��=�`7}k���p�P%�=<�ȕ�{�Rn4��|L�$���gMX���h�`(P?����-���G2�{iG��R�?���/��쎥���4�z�_��~(a�%%xCh�`MIG�,�7���B��.�"^s��h�w/�[��4�e�~s�Ɩ"�>�5p���7����kヮ];A�IF��!�`��3�񺒭dT�F'Y�2>����SV��Ǐ�ێ�t+�R#�k˛ƍI�����7�xc5*(���|����ONĊ2%��%��ȿ���K�c���e�SY���rT���\�U������V����"�[_�FӱZKY�g:qhs�+P8�G�
����Qb0�5dP���2�C��Q�z����&���|�ٶ�~s��iw-Xd.���Cp�B��k�y��Wg�z����A����T��3��+F0<��E���3�=�=�"U���� �(6����d��g�>5E���t\� m���;2v���"@* ���I�1��4�	��U�?�Y�˨�G�����*@���a��%*�O!��v�U(`I� і7kh���v�T:�ٖ�g�u|k���l�\,�3c&��x[Hh+_Ur��|������������H�L?#�3�5����mc=
�o�!{���Y3�/*�GN�l���	.��=|aKC�5O�kd#]~��6h������NjD ,-F[}ܪ=*�V�I�A�Y~�]�ۡ��6Ho�@)ϊJ�e#ms����w��є�̖�ϽiM~u_�7�Q�f�C�s
Bd�G�J��̳�1 g�q�wO��湠���_}��6�\�ffY����ؾ��h�/�Xgě����E��,]ZPp�-�@�� BmF>�%c$�j����ѵ_h��dC( �}���v�(g<]��K@<HZC�]뫵uTmP��NI0#V��D�5����7�ۊLTȝ[$��ɜǀ��
iO��%�^� ��oղ�0������.��h�%�'�g�Ɗ� i���~�Y�!�k���7;��� 
 ����Av�c��
�8���N��ϺcE:���ϻ���1ό[I�K���:#i,����My��p�v���2T�Yß��o)1	A��aF�������x<�q��(kU�7D�V	� �M��:��D�^w#�0(r���O�,���j@�
��0+�����
 |��i���p��f�-�E��J��Mɍ��K0j���C��~f<csb~,��xDŤw��1%gp����gd��c���y��]P�2tg|��b���ț�� Y�S��8�<i��M�(��]��x���.� �ŌO\�w:��AO�� �?���h�2�c��w�wu�H�W��3�Tέ��{�] n���rݿ�a	�O��*�~i����|9�>B�#�La�z>>Hr�!�q�oܛj	4|�|����sv�d���#�������J�@́�����;ekm��2@Bu<FK��.إs!��E3����@~3v�~��A%�0@�G��#n�(4�k1H�*�W�Q'@G�yP,&�ghj��3 �W'y,���2����Qa�MĻ^�ѕ�d�F�����2��a0H���#�Z���}w��Q�ڋ�i���e��n����p��砀R[twl�O�xf�մ151������/����e���6��d��,��T�>,Z����{A�}�?o7L4�S����� ��u���Vgu�����z)񹒳#�
��$��Ǩ�mFM��ۨT3��1��o���r*B`�ǩ��l�9� ��!O����b[=�\;�(&v2݉^)�-</�"�e1�E\(��}����S�&O���E��)�\��m�B�  ac�u�bC����7`��Lb�)\�=#ǣ��81\W������� 3:f�Z^9�cw�[���� ������6,'8��+-��r��
��pQ>**�����
7��,�+�kw�w*/��G�K�` ��"O�Z�zP�$	cq��V���x��d`
�]����]Rfa��LE!Pt=x����Z�/��s��-CI�
n$$�B�� �h,ù>n�u���z�ºJ���	 �v"�!�~6LU��^�͊�%��Z��K_ *T=��b$/x0�0�?�>Kќ����B �M'�T`H����j�SnL��8Hl3_�>�m��7��t
;�a�AdK��}��&�z���C����r��n�Ҝ��{q$��9� �+���\|�
c��ٗ���`�^mG���<ި��"z���Y����N�%�\����>���o�!��?�pZ7�`�ô��wJjn���ܻ�9�UL�X�R��YR�_��:���Pٖ|y ��t}�i������F�xC�����q�'�C�Ca���5|�O��Z ;K<Q9^(1�����T��W��y� +3�e���t���!�1n<�W��Lu��v�!zwl˨���2�����Wq�z��F���3ޙ�� �s�,$f���+ ��(��oj����y�W�	�.��Y���#xw�Q����1�  O�C�;u��tl�(�󭻘�9�co��e�j�T��y��1�	zH5#,��ɡ0�IF|�s�͖�ɗQ^�����r���n��@����o0�j/Rf���;Zb��l�c�|vm�tc`�P\/Ā��]� ��!Ts�\�'A1�� �(�x�S�� n�ѓ�1�?�5�0z/叝�����|���a�X���d����L��f|c�z���8}��������3�ȗ0xL3^�"�m�$�c9F�=�<2
^��5D�eay�I١-�t|M���v���q�Co�z���շ_}�������_��_����o�Ҿ��+G������F���]Z�>5䁕�����__���չ&iԯ}`=O0
��J�7�w>v��|U~�0��P%�g{F�Os�xGK�D������ݮIQst�=�]lί,?�28�e�ш�F�O�v_,<�-N:�̰"5���[��^m����C��aO�۶�a���N���A�5T9rW�-϶���}�6z�®X\ά_�x�Q@uqĽ;����9����E~�3v�J�OB&�� BnYYF�h�R��r�|z	�E@��_g�i��-#?R~p�O��M��o���Z�0��@�ь� F]�	�����6��%$����~0��O��Ԩg��*��{)�1��3UF-u���»:��L��	j�iIl���~�HI�����v��K��� � <����u�L{8��W0��q>�	��a��!�'�D�#҂*��@�,O�v���9��z ?F���e�'V�
��p]֯�?G��,�\���������ǹ�'0��a�q��6�������x%0o)ݺ4��S��t�M2o)���=T�O��G�+��zĸ'˳ꍨ!!e�0�cN���Ӿ���*�J���)#�-bu�ܢ԰���O�\���T8�ed����h'c��i�>��v&��;�T�j�+�k^�����[C?�%F�/eK� C�tU�w�BdBY~����+���4�YC25~^s1�
_�T��i��1ة �efh�?9OO��z�u�%��|�?��nO8��"�ax��.U1��y#YG�ͱ�������R��XF�G/T��H�ϕ��~;�~�$�1�iL�Yܕ�u�X@�g���ZUG��eU'M��? go�o?8��t+v��E�@b���(j��ä�'�.�<Nh����3��gB]���	=�>���}���U�Y�U2������|�)����^4���{��Vo����VVgq�FvD�t��O�:�T`*�&X�G��ʱr��0��LO;U�>I k�Xl��ʕ� ���]pWb���$�ID���Iv�i�h7�C7�U�"�p6�q�w�U�S��Y��F7~�"g���4�rgUݵ1��%j����C��1�y�����9������39��@z�b���|4�Ǘ>��er�G7~��� -���<��q�9|P�kݎ��Oһ�:�{�ʮ���#���B�V��3��/SaǈbdiA�)1z�B�&ܔ��V�6�{��o�d'*���F�&�7b:0�ڦ���akW����F*<�ꋿp�j����6l��ZL����(_�3$�ߩpZ��q,?hߓ��KH^o4\��IY�n�$Ͽ�ɃG�0r ��8+ݎ��uv�?�+��o�h�\�R �_K#�N�-7���"�^��k��L鉹����e��>VР�0g���Y~�)7ZJ`�
��<K�|(����Ȗ��퓻�\�b��d$��ػ��s�m������1h� �T3�F��y��k2�,m䫹ſ8c��r�ȷ���i\��j7 Օ$���n��B�D�[0�s'oIVC�IDH���
���7n�į�ni���շА�K\Bn�E���Z���b"�8����[���[�A�/	�V��;`�U�������ḱt����'Y�b�\w�f(����1m�i&��ލ�(����!�dH몥�[~��	��[C0�*Վ��A��pȚ{7j�<x:��(HHu4'�[fP�~Lz���P0v@;"�2��G�4ǽ��цG-�~�j��F�z���.�ye%�]%�_D-�F�7_�ʸE��d̶j6]�@2*�O{lh��y�\�N�ҝ��R7Z��ep���xu��(�t��e54���@�UK�2A��1����]�	�y���o�^�*��D����9	F�Wj�Ѩ����W���Q�D��T�	��	��8)W� ���;�6�6�
0r��lK��s l�ү���`�x�Mo+��,;��,�ӊ���w��)��]��F|��]�g9�C�+k�J�8�B�jA�Va(c�^`t��>9�5'
(9_}R�|2z�tX�o�Nk�- ����ֽ��{ҧl �`u����ͬۡ.G�^�eȻ�6W����O���7Q .qK��Qi���e���b1�Ϊ�㣖A���������k��I�G��R�I��f�>�l䀉/b[�cG���b�C��O�����}c�]��B�����1y�BW��4��a��~�6';���տ�V%��EMk������pR מ��4�F}�q�v��������/]m|9��55��YD2͎��$IF��������2�Y�VB������n+�%�ro4̑2����)}u%B�"�`���a�P�����mkX�Aއ2�:o}�������@������6e�ŧ�ڻjX��Q��v��ZH�l鮗|'�Y���)79��5|�~RN�%�7����e��Q4���eTȁ�n��F)9��h���!{��^�i>��FE��&w���G���mW�u����R���қ�U�6�v̐�����7Fv cO��M�H&��+c�fA�#���~�J��T���P��ڌ��Q�<�i��1�L
?�u��A�(%��^_����$�q�z���[��&�c�`"�e{�=dp�a
"WZ���z �[H�ߞ=�O��ظN�\v?>��d��<�٩ۏ���#��N�;� �P�:�H!D{�$�Y�HT8JO���	�8�j04�Le^��E�J�<X�c�R�$���޳y5� e�sh�����you;�|��'nr+����;���q�9䭪�<��1��Z�9��a� ��>i��#\�˔��`DR3��&977j@tҫ�k#�*��fk�ֳ�s�_�Go|٫$-h\LwT�	p�yX�{By���v�M��BVw�.�k�� �������_��y=4������u���%������ߊ@�H<^5(�o�2�0��՞�)�ҋa]Y�j�u �&َ����$$�4�Ƨ��[�0	��_&��`hq�xr�M#�z���uO�(��2>=W���U��J����^�<�>B�N`�aV�����W}ѻ]n$4�GG�|.l|��8�s?f���럚eT���SO(US�,Oc����2�FƁ��@��0(��d�ضn���v���u+��B;Y�XQ��	���_��!�!������g� �)����7��<�W���P�h��(�4�<ډ��hz�F7���=�D��eKRӄ�.^&�C��򋻋N��`��矚Qg��*'���׌�1�%��*-�Z�ږ��J��'9���-�1���v���:P֨�:XY�=@CXS�xC4��d�}���1� Ð�����+ulA�Y��J��hEQ2AZYv���l�Id�䞨jF�+ǻ�!#�~)� �ƛ�<M��zK"#�X�2ΠM�t���@�ȣ�Bj*3 ͜�(��p��a�2B_�R\]j�;p&����䟠8r��1MU�?�p��m�dB��)�G0�rn��ܖ��C���C���č�v>9;���v���(�~����٪V9*vE'�D�Q��z ׁ@/4x�B�[���ض��q�@h A����{�Te'Nv�Y5�jΧw�T�A$�q��0��(ޮ�%�3�����+'���b�;n~=�q��$�Ӓ�o�v�[X;rs����E,�Ez,Y��5n����_�|�9J�܄�L��KI�ƍ��HWn�o�U��+��r<���2,!��W:��?�~�d���d�_�jF#��C�� ��B�L�cY�,h�H�������Sɘ�paK9��J�t0��Q,O����]�B����T�|�AېQ�����Sc�)&�:(�{��M��3�!�1*Ȇ�!Z�=�hD��L��gO:���X9[�kS>�Z��XZe>�l�q�l������fR
I_��Q�,N�ș�}y�h4�27>���r�Ʃ|�i�!�Uw�o
jY�@� ��,&��+J>�{)�k�j��xH��Z�ԆN�ذ=�n��!1��˛�Ι؇WJ���ُtw�_qn~�*8X^R�='OXk�0R��>��9���L5��gr�m��d��qzϩS���5Z6�_H���Ĳ�S짙�Tu�z������`BV5�}�tsD�\���Ǩ��o�+�ygl��*�+'#���x�Ǭ��{�|zW��B�ܵ�/3��No\��8�m�\��j5cD1�����f��8y��GhPE��SǗ�Aɘ�~B��͵D��B� ��޴,� 5$&��Q�����֩Ҫ�R����/'@:T�)@N�sc��Z�Sc��-���d-�𙇘0s���c�6ɼ�WS�ސ�÷��Jaȩ�"4�����~�iT������2�G�8W��}�6\�n��}���������r�����t5�Yn���6�F����V�e�VR����`��fRh:�F���1�dxEԓ�f$3yp?kN�n���@SJs�<o���@�����u ٹd��[��WԻ�Q���T�a�P�N1:�u:��t(BT�~gkO�#~����&�2:�XF��Z�Q�����s�o<qaV��#�[�{XtT�<o]��p����⩛x�'���m��<�V�C4��e
)� Ħ��h?=���K��@�$��V��]!�������W���|(@^aR@x>�����%��񫔍�����(����{Y�AW��c��@�	�7 � ���]�a2в����k��-�N�a;����T�5'o�=�9�b�f;�קE%6Fp-��$��]��^O�=kQbֿ�S�������!F�Mû?�Q}���|*���⳨��oW^�(���I�_�w�����V��OƊ����v!�ш���U�9��n+�?���õh�vj�(��=��O_em���Gj�c��/�����܊�(5�zܨ�(�����9/A
�+&�~��w����jK��B-X��Nc��:�W��?�~��"B񄳀db.yi!��coՄ�)@�bp�ċ��ikM��&`9�
�g�͑{J^�'����GG�b+b�w��b���~?�(�E�MY���͓�lm��,������������g�n��NG����^f\���<�#��'��/���J}����礶��+��
�D�,��;qP��rُ�K��'��q�f���	�����ۭ�h�,�Tk;(J�1_��>��U�:n��K���HnH�ZIn�<y�Q Ej�(\F�_�cm��x!����1H�}�n�l�w�7\��n��;��&g������C��8-�[/R�����c\-�p�>��VW�ۡ�[)�hۙ5"�<��JRc}<�R%�B�Pb�~_I��l�Ju 7���LB��4����R�#��T��<f0(I�j�z+��Oj�)�Sm\&������ 9�a;l�H��a�h"�h�l6A�1�$�G¥h�C'�Zw�1J�/Ny�^fZ�es����Wݿ{w�Ġd^��9���ݠ2(á�����;f���Z��C���D����������a%���_M6���%�}��`ղ� *��4�ί7^Q�)j�2� &C.w9���t�F_���J�:��
����k�����bEcs^B�v
5�{<��t�mii��z���?�{�+)nF�7�o�m|T�m���^�𵝴�0�XcZnbe��Q����+D1�AMh	%�
k1���{�˨Tz���rg��<�I<*��)���*g7~�x���<L*���Z�+۔�ڤfU��vSӑ"D1iŊ��;m�3~�W�ӛ!F��~�_��}�\��j=�D����{ݪh,C��蟋]�"xx��}^��#�,�?̵GCNiI��q9QF���uy	]�i��P/55q�O���}�h^U�HXr����c;y�Ս	�4�8�Sw$a>ۂ�ɻ�b@�����?�7'3���AԴ��oǊ����r�Q3>dQ���F����T������lȘ#*z��'� +�J����y���7M�0����-�X9rĠEO�+7����$�����DE'C\ifb4�բG4�w�=}nϕB���>Մ�����^�C��[9�!943
/D�6����r�$����2c"uk�6�<}fv��	
��jX"։�Z{�=lH�9/7 �|H�E�UA��U\��� UjÃW�Ki?n��P��Z�����+f��ԆxN�K����	x/2E,���|��̉�v�о�,v��6+}Fj���4�]t�s�{u�Ǝ8�+�r��`���N4�k���(4}<~=���5k�}f20tjǓ��q�]���c�dyD�N��;r��/M�L0�}?(!`>��1j?�
̉!8/�G�p:˝o��v��U�A?�3"��x�!�(�)�ۊֶ"� ��[�0eg�_���-���R9,�"p�X� ®��͍���y����oW��؏Yڲ��?��+�5���@���;��l{�R�y���8���,@��0��@B�;-��_��b(��J�'������;�����J/�ڔ�#ϻ]�}��b�͛6������~� v���Tҗv�':/ X��֭l����;��n�1P����>PX��UMj�%lK%�%��.@�H����"ۜoDxF=��a/�
����tNT9�ݺI�E�?�t[��aɬ���R.Ʊ8��s}}���k.�>`���>wdW/��M��H�̹��V㎅�4��
	�,��Qv>j�M/������e�����ix%��uy���ǎW锂
ĸN�CD��R����{�O�P��H7=/7���O>���&�֨�+*
��{�4��iQo��b9@�4'��Z|�4{�H��iv�������A�n����>i�v�Q�y��({0��t�3B`����A��x�	�G�8��N,�$ �@Zb�!F<X^�O%���ԍ̄\�>X�����W��ʬݼ���L�u�g~k�|��3�
�S1s@h�\2?����)���cU:�^yy��lA���dV�kj��<zs����x�I���,#�@'�(�f�hF����L���p�79E��k���@���?��lF��d�z�a7^�5�F�fB�n�I+R��ҭWn����z���hi�F ����
�?�D��~.�g=����}n�ԅ�fۮ�
��)�EkN�Wo:��آ��o��ȑ���Xh?�U N�XӬ,O6c�=>�&b��,=W���{�T��#E��:��5���˰�&*�jxP��:0�g��%��2�ޗ�S3"̰�\�|���#I@m�)�;F(��83#�b��Z�-�G7aLF�XV:���)��v�ތL[�<D�c7���^����<{-�-�{����S���Ճ�@�I��sxfƘP�
�2KHmf�&u2;��)C_��-���#ݶu�o��?��Kvy�=(>Ɠ�-u 傕�]Ξr�3o4��]�hL?�n�ퟕaP?�{5�Y}�9�߲v#��/����g�٫�qO��E�x%�_Ց�����B�]Uv�����t������;3|*ŏ�樑�G��9d�O/�_��ͭ_��=�LBdd�Z�k'��9�լ�\�9�ň��w@���r�c
̙����+U����IFw��K�v�v^�����
v��5t���/~p��_j\I�75���&����`�D����2:����\8� �u8M5�nB��Ix8|�Y���P�I���ثw�d�E��E:l���Ϸ^�P^�h��φl>A�[ ˛O
Pc���0�������Wڑd[���^�ɨY�K1\�����0�Hm_;*�=��Ԉ���U�v��OO��
G��ː^9�̐\w�ۮv��y�NUp&�A����Qu���Ʒ��������UB�lK�u���#=`�#4���95��e8�|3~'v'5�x_�|)� qUv}��^��qQ/��#�je��g��ވ�@����bJ�5b_�-�FS'���3$v"Gr�nq��ה�R�����xL�*!8'��v���^��A(��'M�"y�\C�k��"��RVc�,5�x��4X�[W�^�q~j�� :�=(�nG���>ܴuu�z���l!y�lH���Gi��_ /R��*���'���uU�%�4P1��T%Tu �m���Y��73&i������<��)R�2Q>[ֲ?�W�坨��4�G�S�芖8�[ci�7�=}g�</O�Y�;7�u��U��q4�鲼���33�G������vo�8��Q}��$5|0�}�:!�G���>�lg�^<64c���A�m�)Y�	od�x�U(Tй���ѥ��䫒I�Ɗ����/w*�d(�U�~��K��>�K?)-8�Xj��P����9^���YyDsc,7GwEy�+Ɲ��9��\��� O!x�0�^�����D��@F����l�o���\�̃���6O0�F4i_:^%W��n�X�#��>9�~*SG"�XƸQ��ah�Ȅ�7G=�'7�L��9)��Ș�ЦM+G�E=��ba��Y&�mΧ��I�Lo��Z������iֻ��l�!�i:��{��$;�A��G��a�H�lMZ]	~Ӎ���bk.,%ͤ��/r>^��qܕ1�=�GW��|�B�u�n��#���zEmR%Z��B\(���rN�R�����ϗ5ͩ��_=��U�� �8�'m��h=������̫#�z���Db�D��8T rb���j�K����N?![?���b��Rh4�O?o�Tdq?�h��P(�V�ԍ����ʡ}�N�w�h0b!�>�DMG�����A2�Llc�iE�[tz׈��;��\����u���"�i<*��.j�����Բx�wV~��	���5K���x�BظG�yy�2ݨE:�'jST�H�ۃȖQ�鰶b՟o�P�,f5�:���>�n�Y���~+r]=S:����!���a���������T��F��3ٍ��g,��o*::�o�3b8�+�\�͈2���'!)嘒,op�b�	�Ǖ�O6 ������.g�Pm�*h��?~�4�y�hc׬2(T�|ҀUΗEkY-� 9���?�Ċ�[�(�1^m\ Hᮭ�cVS�oZ�~�`398�A��{�v��z�#']�8���'(a��Z�f�S�P�Tw��D/���t[��kǽ�ń4(�+4rH������j$�+UU�Zb���'m����m��)E�3_!�l&�s��=A������;��'�; $}�Z�����9C ����+�@qI�=�+u[�M�.���x�2�T�L�7�D�o������¨�^?mVW٫���(���I�$d��E�w#�k0�����Z����V�T��1?������Bڰۑ�]�!���;Z��n���������oj��+U��۠_���WPai=V=�kXDz�|��!��H��3!;�"�<�*����2H�J� ��o��w��P�~�oj�R"�֭� sj�ߧ4���?B$�?��L� Q�ո�Ο
HR�~�iu�˯^b8��S���$�+k�
43�.�6am|1�6��Dy�[�Am{�*�WF`�MT\ft1��J�!�{���	�q�i���O!K]P����4�<1Z� 	(%= ��"27�%�M�"%&�S��p������s�ܑ��1B1O-��KKTk9�~���Klc���LU!̧/Y�o�퍍�P�+��Q%#ϛ�NVU�\�pG��$4���v����r.m�f�Ԕ��[�KoO�7�U=�h��8��*J�����*�F#ga;>��x��^�Ч!1W�{'8xZ��J�g��l�tzg2�14R��(!6e*�٨w�����h����Uey�����j��3.�2GПԚ�3։/XVK'ͯZ��sٛ�l�f�k��,sE3��F����٠�|{��|�[�c��
�d��y<�pr���d.����x�|X��;��GΤ6F�v�p�,X<��l�A�5��/�/0���Yo�JWV
z��8n^�}�ǜ�ңۅ�!�z>��͸sT�y^]��j�"[2I3�䤦.Cd^��{*�lvȇ�A>�0'�=�L�>G$,�'VD����pԷ~�iT��-De�^uZ��}C�k�\��QG"͘��q�{S��5��O�h�D.s�*�n�,qI�u�&�9@�PIq���S'�l�^��`=͂�B(�Ca҂���=(?raOB�}�`��WH���Ygd�%K^��X=b�]�}�^��гzT�R��D7���M��+�O^��Z�-��h�D�uܝ�P��V��iY�� �}�e|l�U�5,����B�����$+�z��aί�I���k��{f�Y#�r�a����]��d2�$K�QR}�C���Ɯ$�ht'�g��8L�����b�J{�U����KDft=71쨵e�F�"���ԥ�{�)W-ԽS����-�P�ɼ7�Z0��XX,l�癬��}e�7��5_%��28[M�^1�H��@UU��i���2 ����21>��Ȉc����fh��)	{q̯��@�~���E�rZQ��^�Ȧ�}Y��*�v�4�����%���R�#-�I/�Q:��;�lS�n;}����%�k��W.{�c�7}?n�Z�;��'�q�N��#?�����5R��{~�~m�� k�I��[py�_�O��uK}���Qj�.t�ￗ�pZ�S���-���B��/��B��/��B��������oRRߒ� ���B������S�J��
1�.����ߌ��v���p�c�OJi���no����5Z���.5Գ(_<�>�V�xO3rc��`žK���酱��^���>��b��ӧR��㗖�II]�i1�zG�(R)��MMbo������B��/��B��nΉ
&�#K��=�I!ӛM���������Fj~~��y�*�P��V�pc��=�_d��vg��#�S���ۤj?������x�tU�[vm`�z�\�h�)^�9p������K�Z��2!y�I2�g�e%s��yL2�%ɜ/>����_|!���_|!����fCOwJ}��ڴ�e���k|+�f�z������x!c�t#������w֝mj|\�,�,��������K��PK   ���X~��k�6 4 /   images/663b53f5-e86a-4272-a51e-f5b809259b46.png�yTS��6D��U0�*�n�4JTP��� ݠТ�
A	CP�y��j��mQ�L�4�@ ����@E� 4$"B� ���пw}�ߟ�ֻ����^<U�k�g?��u��/������[��O$'nE%���W��o��� ~,=󟟏|F�W>𿿦�t����G�ɩ#��/ׇڸ����;�7:D;s���(��_��b�	�3��G"2G))�)	�-�H��[_Ɨ�e|_Ɨ�e|_Ɨ�e|_Ɨ��H�<�/p�������/���2��/���2��/���2��/����bl�9�Ϸ �?��7��S�9gζ���Mт��řv�����'�6~�t�y뽇N�ugKZ����������E?�G�'���O�0^}b�r/��̪�=9�����g4K�?E�d06:�b՚*������2��/���2��/����6�!7������CSoo�Q�ا>�:��3�"�ܾ�yT�_Ƴ��1\�yk8�v~�V�����g���d)N�.�х�I�3L&�}z��U�B����I����Os���:�O�@�bt����j�A��,��YZ�Qr�p��`���5��^Jt�l��3g��g0�������ҀŌ��~~�hcG����a{	|�K� ZZ��,��%�o17�����2`�`�~r�p�*3�������(�w�2"Ɂ���@�hy��ON�����x�*���/lU��b���].�?W�-�H$+
?����%{�1��x�EF��*�2��K����AZ�� ߸�����4@��_0+��r�� ���g��O���D����N�ʲ��\�C����6t2*�vnȺ_`�",������Y�;����Ui-j����L72{=��H�5����CB�:�F;���k*�3{vaa�q5���[X@���n�2T7Nah���-$NTײ�ڐ�����	]�8�scO�*�XwF��)(7�x��xλ��r�	�F��(��s�����1�QP�Ƞ~���4*��M<7p�'��Q�A�����"�t�A���t���#ڇ����l4}����c�v����b�|bTx��DǑ=���M&BI�$������.�k��>Ը|�B���C��VQ	Z���L:gO�]9����C'�K�Q�x��ߵ?^˫�S��ai6Ǘj��:ٗ�`4|x��Ǐ�_�~��*Z�&c'ո����L.����\쓷RE���a���<�g�$ݽ��̈�r�3'�0J�����:=�3#��a+�^�V��65�Lm4�����Ne��w�7S3�9�70^0�͈����Y��K(��34=A�)WB�ێ����%`	c�y��j^�1��!���Rc�	1�'��p�<�M[`L ~��*3���gϞ�~zi�����'��&�\f�1#��4�j����]IG���C�������<^ֹn̎�1;�CvOm4��bD������:����xY9_"�ğ{t{[!��9�	�9�^��I�s7��'�b<IT��V��1 �y��lb�H
�O��ƞٍ�݄(�S@���<H����$��Q���������*�� jA2�Zf9X_c��i/Gӵ�����={6(���������	�#���Tr{��@y�?~�O>����~c/o����J\��ê�Ȼ��sQ�T�&��`j�11�<�C��,��
NW�M��}�*��<�~UhNHLө�����N/M|z�u�~zԳ@��}�<9����>b�F4����eЈ��Ӎ��֧6��0��D�z���j�4 'O��
TL&^rd��z�s��?�iV�c���4˼��i�����^�� w,>�qt=��c�H�����¦�F�������To�z�b�!~ԅN�m��m���NAn�>13��wSEB���H�zE�^`M��F����W +6fo��I(ƽñ�5�!L�~q�"�qP�ܞ̜��g�A��m��+*��-��f����-t�3�B�u�9��`����5����h������;�s�F�,���Ը���3��G_LY�f6 |G�����#��n#�[K�Dp6�x��}�o�=�{��x=��b��r8�r'6�̉������.�\��]��wz�;Ñ��fG��l������mG��C6�$�'��]���drd��ߘ�F�/�M&&�3�/|N�^���7xօP=\�ۭ�
2�hƩ�VS%�w��>t7�ޓ�lu�;���+Qm�YP�����D7y�s^N+/����{G_�\��F����x�|vv6���	e������?lf�J�����ߧ3���_��- �:�~>�fE�Bp�:�|G7ӬEIĕ�@s�&9��ͼ
Q33҃t�b�\v��=��7f��Q�n�C~��^��ӯ`K����4d|c�3�p���2�����|+3���MhN�+v�՝==D恾_��.6��3p	��w�t��(�EE �B V`��Z������-_8��w4ՓL�VJ��gLSɱ�eq�.E/�v.Ϊӛ`j��������]���	A�u�ݾW�jS}RwCu]7/���E##v##��-���x�'w��}M�������r�E|+��Ң�����A�@Ɋ\�Ew�{��]G�p���̙d�a�t��,m�_Ѵ�����������_w�F/�PW0���Idjw/�/��0_:���}��9)�s�
?t���qt:�SS`U�jh�����]��?�ÀBj:�'��/0�����q�<쌮7'Zs��u/�jF�>�U�,�T�;�O��E�t"�qF���o0s(G�FzQ���jpئ�sY�c��'�A��)fNkK*�}���ݶ���ej�W���p:0�
n�I��,��،`T�QR��W^^�>5�9���=��*��U�쩔��mD� �y��z�E)�lA��i��v07��r�m+������X4�;� ��?�ɖZ��הhiSS��%�%X�C,���:\QΏ�$,���.������?�.*�*~XW'�KVw�1���s��C�J���|ud3���F9��{��̈�EZ��B9�If����O���0�O��K�B�W��6Y/�>��X�[���]X�|a�{����x{ژ��~-��b����@W-��z6��
a׾b7A��=m ��g�26����6�K	�bq�H�	D�	��6�dE��=���f��0��܍�!뺺�ɽ�F�������_��Ved�%��<��陙>��"
0v�:b�(Z� �F�����cG 2T�ysA��0-�Z֙�O�U�Db��L]��,�Ί�֫�����J���+B��&��>�e�Y�X����<��s��y�,����r3T����H��ŵ-�ڋ����y���ڨ�eO�Cql��G�a�/cz�f�l������~�����ݻwS�b��,d��n���0Am�:�R 1���L�".?Ƣ����w�j��橐�]������+d��b/�S��E�JlA&R=F]8M*�.�Y?=�}~W��ѣ3��l�t��[ I:_��,���S�NBG��S���Y���"��o�E/ߙ�eJ&��#�1�% �0�t%C��y�n� �G�Z�="��K���LФ����?���;�`:H���pc(J��)�`��bL��ئ�ZW�c(G��`%驲v��j.ڵ��������B��@>���k���\�7�,�h��յA��{\56P�O@Z�'��!�Ȭ�@r{��H
ڷ�K)�!�L�� �;d�f�i#u�M��y?���A-���,���W!��x ��Y��ߤ"Ux[�'(̌�y��Wi�L�DD�u"##�o�R����N���"��&�����?�ݎF�"��p�U�6�E���"%���u�s{}�C��oѳ�A�����踙�7�C8�VO&B=Ȗk�Ҭ��o2�3Jk)�m�k!(�̒Tn��h=K��L�6a�X��Dn��)参��9}���Hr�2�b#"h#���
���Y�bՁ�G�g�uT"���+��Z��U� ?7rX4y������<�vP����u��$�F�ҙ�.�71��
JH����}9 #6�'�@'�tHc�B��Ħ�>:@��xB@��fjY�?A؁��M�ΉN�aY"6W����1N�����=t�����{�Cn4d'Q^���Rۋ�b����Ug�ꔵ����������[�V~���s�1���Z���⩑�S~���'ZZ��+�TFo��O;�pZK�J�$q��Q����U�j�0Ys�I���D�\*sfpp|Z�p�Q��%5Һ�3n���?�Ŝ��{�����n�1;�T���0,Tl�Į���.��oMd��%Q`���ۉ
��빯Gd�FL���=�O��+D������C�y�`��>���D���M65�&ƠV�3��_&g�2����E����A~q�_��j}ʹ�vR(�ܿFP~f�U7w��G��%ݩ�w���J�2]�z��`���-TN�-^=�葆�R��Ϯ�K�7:5Ǧ�58v2/f������\w[f���vl ժ�?+ ��M��U_a��@�y��TF]P�J}��</�o�d�(b�'��Ю�yi��k����t�RI���<x@�bo�w4R�i�z@���t/L,�l��Ż�E��9��#�P$̔�r�����n��D;}6z�:�aC]��r����^�� �ÿ3��:GA���������0p4�A����/>�=OKcv��'Y��>=G��:'XO�}܅y���k02^�-�>�T:�z����~4RN��蚾=�=�x���\��s�����4����ⲟ�u�\kc��e�X��&L�a�_ �[�sl<M�u�yٓ�,�S\��Y�41ܪpk�	ޖ(j�������"ń��>��xG(S<��]$��s���T�؄���o��?���~sÃ�#��= ��E�@�����Қ��b��Ӝtz!b����t!�N����ǟE�ȟNv��������� ��.���ZW]z" 5Z�~i��co��5�b���ͫ�q�y�[	����R���%F�b.�|	9��k/�&.����������Q
�ѧ?1��g}䝍�&̘(R�-i�s����5��W���'���X<��1x��_��'DNM@��tu�u��#�W��a	��������P�34އ�`�'��R��I��!�ꆔ��쓁��t�jl$���"6_k��xqRV`6���l�p��Ю+ Qe� tW˿yr���!�/���'5��c�ׂ�4J� �S��G��#��7�D͑�>���`]o=�,�t�9��=R&�MC/ӭ÷k�rѓglb�jV�Ps7��t��1��rF����A�%\��9:�}����g.>ygo��E���|����n��ٟ�~�QP�4,`	y��7)b�[Jpq���1>��V��,+��w�^�l[�e��,�U!�4�p��l�쪍y�-^y{�9oP�E�f�o���*����͆���|���^���X$�^�e������`M�K�x|,���s�}�Y�T�Z|�~��_.�)�j�̴bī1�E�
zvG������`�\�t���Fz��s6��0b��5��9���~�_o���	���?�h�K��T���k����կ��śĀ`BZ���Ț"��wQl[x���	gM~�T��&�͗�6��[+�	}��&�Հa����0�K��=PP*��0^z�n?����S(���1So5S�Y��E���˜I	��avS蒶��ܓ�/<D�����#�eޙ��
M6$�m'�c��݋9�gw�e^ڧ�:5ma��o������b~v�C�{�W}}����JK�UY�
�Jc�yccc����<U���E���9YL��Ւ���wA�e����Ë=�E�����*	��XY2P) ��-��t)8aKj����ж�*�vk�dS��XZ�@�x�SSr����D��Z���,�x�M�}*;�0p��iqjʥ��o�y1� ��G$#��N�d�zK�2�}(��?�|�u�V9�'A��1B�nG6���kD��c[ݎ��Ps#i�b� W ��->M�,?�'�!�� j�a�[�`�8� B�8��W�/j6��%�C���b���mܟ�:�B{�����������MaA��Cq	�k�
���&h(%p��a��AXR��~dM&�h��uR�������,sٻE�H:
��GDߛ*g:�	�_��[7�&1l��u]�W�2&�MXo�u [ �p����d�Y�C�d>��w2����@+(��T�2�#�@ �)cF�#,0 �^�K���5�j�D"����;U��� Egȏh��}��B�t%}����G��27"�0�(���I%�:�8wGd�fUUպ?���6�8�Js�
��)���-�@�ʟ�G�ز&�~T�C3��^��suc�4�]�ɖ�Ѥ{�"@|3��Q�&�~^o�l����x��%D#Gag��n'�@P
#���u
����b� ?���(���13�~K������6LH^�o���"�Vh��c��?����#5�QNiڧ�NM��JwJ��Z�#�񿃏�7��𨋙����.� �l�=�")ox­�$s�����4�Q�t�0����c(��dJuT/�tCI�Z�kP����my���E7����zz�kC��߀~3��>t�ҩI�� ĸ����T{�z$~�*�z���4ˡ��?�٩�,�w���h�m��B
�����g��]Cc�YT#,�f�L����"�<\b�h�͟�+�5MihWTG�am���E�i���a�B�O:	�˹��y?�dc�a�"�Ƙ�,�����&���d
�Ks�i�@��v!��6�Pq!9T��3�U�U�Y��j���L��2�o�1�ڊ�[z@��������S������lz怒���y�!����������#�v��)�A7��ߓl��[�;=��Dy�d�`����@�W�|�!��a%�H��+ȉ�m�'t��1��0�	4��E�^���l���#̾�ݖ#���yaA+]�ۿ���O����a˶�㫀�ܹ�Ҕ�P���7�U��U�����P6�#w��'J�kC7�a|�Z��XS��A�	:�'�9�*'^<31,��;�NV��2#� t��;O���QpA��%q�'2��<g@�b��G/˴uu�� �]Z<�������
�=|��`]W���l]|{�E�	�V�d+��Uw�r��x6�-��h�����*uтj�j\O4�ßMrjrFHJXr�xX�F<�A`K�P�x����ȯ����T,_��Xm�N
Z�Dr�o릱����cݘk�%��E ��:�fek���N\$ ��ҋ{+2^(kݘڨ����	j&�\_t�vJ�Q�@ģ�v�z	Q�$�
�}�Oj*C@�pC�`Ț�'�{��k:<��q��&�$����;�����޽�c��S�T.dB�2�`�����o(ZR5�Ӈ��ݮ:�H$���X�y����j�T��wj
����.徙}���kTAY��TU8����WKKK�� ֗�|9.��t�ZR�e���D j䥁�2ѩ���8�{��p��I��kv� g{�`�l�%H� ���NfjѠq�:�s��]�{m����p�3�����N;��*�%�����1��;[4zT\fJ&��re<����^܍�CB�5t?����.]r���BI8H�i�4�P�W�(�|�3�`���N]��� !�v����q��<
�?����QX��k�G)�M����ԖO���c�K�k������I.FU��=�YG_��kD���k��n�����
�ljh��&dHۛ�#
��֎m�rA�Am�`~�a`&/�$����bs�����0��˥��6��l�!�1V�� Oͱ̥��#e�����\w��A�1��҈�ҋ�|�����K���_'�E��sCﷀBQ}�\�����I�?k�&/�v��Bv�M��2[R���~mo����z���sf˨L+4ӎ�
�k1�J�hٺ�=]�!�
�Y�����N�ꦢ���0���6�BG�)ׄ6��Kq�& :s��U�#zĝ�țnD��k���{$���}���y:�>,&fn���$b�3�F�T�f6?�������N8^ָ�$B�5(�d��c��g�C�����߂�V��
3'���g�U���O^gm5���@��x��#����_��Pƿ�u`���_	���������Qua�G�0��x�������	� ��)0������{ī�o)9��n]@ݮ�������ӸX21Pm��
H8V:���a��|�ۀSl�)�a��`�
3%�S���'^+�4nq��
W�T%@�m�;7�$#͗`��N`fa1w�C��3�/���%�����P)�झ���	[�]^ܾ���ۋF����ə���t������@����)߿Mw�(g�f{���z��1�~|�H��?�鬈���@���V�܎p�}�?4�3je���^�^��y��pKl%���HΝD��ô�(������myl��2�Uf�sޠSS�Tn#ޜ���>��w%��T���aq�0�P�kk���s�څ[	�91?k�]��Y^��nV��s���Vtm���js{����8�yF����ů�˃������X�����X��E�#f4�Yp���r���\�|��&��/ �S��Ry�~`�R�q���tJVVV&��O��0Ǭ״HGGk����0%�#��VRr�=����$8�mĉ,aW����)�y������W./�/ȁo�`Q�f��,��`&32�	go"�?p�y��V�L`ַ� _8L�rCP��C����U���V�N0����C��D����w��(o�.�l�"rL{[���B��NI�J���"�q�S]�s��G��=�(�yi��7a���B�N�6d�ks�����a����;��C��oa�\<���O��s�7n9!��qV�����P]X:R�)v�����
jY��?˱�@�Mxq]��mp�J� ��L���f�2p7�1\�ূY����tY�OX�@/{
uKEJ��^itgo�v��X����3� ��""t�N9���.���A�~O�p:ل8���(�e| ��h<9�"8��B��M`������CuP~�_���/�����N�֟�V~�}(�KuS����)M�Ť���Ϡo��@�Qx��7�"Vux
j�Cq��uW��x^'�k��l��u���k�l�?��������S L[z�@��;!�]J��)��"E'w�����0x�]��kCE��r�vAX盛�o�?��O P��5���D�p��	a�O�0�9B�� �T��iM�|���[��Wl��5�ƌӉo�D�@���)�խ�	Mt����9�u�E���yi��Ņ��V'>=0���#��!�T�5sZr���������mE���C\���w^�K��x'l%w�t�SS�u�Xf`�~��1E\f���si6�N�G�>jTNT�6��ۧ�po��jGGGb����Adsj"�$z:��{�B��r��>���a<�e�$����p���x��s5����!�9���0m�5�.2�%�z�� Z���Pu��})J��̙x����˰:���W��᥽~ry�_�aY��zJ�"�;dj�i�g��Lk����Tï��A��&۟V�k��=��mi�	�N���;�w�Z��J�sv��ّj�>~�����Y#���{���|j�>�������a�UNv�������q���+�ԸO^���>{�uC�#	�@����N�n���<L��V������e�,����ss�P(�va��֜��'�H�/ Y,����E�/��+�^�v�C�<�mꉹ@2���+]�"��~�KP�5hs�,�/ZlUev�=�����i+�^%�G��}���pa/���Ga�	H��d7S���^�0���d�졉U�v^Vq�`m叫A骏�Щ����(��9g��ʾLf*���R��TH��I$�(��2[��G��:E;�+E��X�O����ɰg,,�����#D��{K��;��B��,�Y4� ����ҴO���R�Tr��a`A��Z	�Kg'\z�^�4�;�,ςb�n��VB5�Q��f�'�0��������^�ϊ��	½��˲r��i*�Z*�s�;
�������U�X��:N�����J.�	�Jm�ވ��E���cK�78�Uw���s*T�*/4B� �_����?`%�׮,���P��o�\���}���G�`~��2} V.�;֠7��~t/��p��f�"�����;v�\~�ͯ���#ĉ�\��;�\~㑮,V�p<b�6ݏU�
v�:��\̮��Y��u�#���Lv�	t�?�</�8lM��aZ,�9��1j,�l�MƁ��cՒS��U`9�H6���|(IP���;*�5��%$��䍃���.���Jl���0`���E����e���!$&8�z^���	O!Z��C:t�=z�(����Ϙ�8�"�`p�����ea+K#�������כ���T&�T�[���L&�771uRyn����+���	����l�p�n�j@#:7�w.�ڝ�K��-����S��4!J�aKH��������?f�1����cR�J�tz�,|�+��lq �l(�W��[�W*NwLaThkiYTayv��d�e_l|���,�ͯ^��ޢ�@�ZW�H7r'K��t7&�/��.}�؍#T��@P�,�С'�Ń6������R�g�d�����u�}������5���.���m�Ɲ�qb^Z
�{0���B��}E!��]�����'��)#�ʷ�^��a�6d��ϗtvuE����<�q�����U�1#��
[���R�u�]��
A:����sNPpp�]Ҍ�0�w�lMq7h%�)J|������w�ޥco*7@7��ߛbq�f�kXCԱ^J��֨Z�o3!�d�)P},,�ſ����x�yԯ�3ն�]˹����]Hk>1��y���9V�8h������a��L�̨�Y����8l�	��Y��oD�K*��P���}���)֟ڮ9�ȘNB���(�N�^i�����7CL����J��$��맢^�4ɟ�Aʤ�*�?���@o�E��/�͊˞<yR��+�ӿ��~G\���������_cƿ�����j��CR��_�`'�k��G�w�<�W*�Y�
���﫽�]��@��?�n��n�0�4�C����Za�e̪��8{�W`� ���/���(ͩ/n��P�b�[�}��k�|-��C��e�c��6H�!�,��Ĳ�^墢H��X(M�%�����MΈGFFV奕�;���=���X�IX��a���6d���;��w#��1[�V��<k+��M�',��{	�v����?�p��U )�@Juφ�:6�
z���huê��| �*(0pޝ�[��{/�ĿW�p3a�N����0�fjj��p�5J���vg�z����k US�Τ�rI�:���ψ*���D���j���+�1�d@\��=��Z�=v]�b+�}�?�k�H+3[_��`(t��ѹC(�ϼ�X������ٻ�{��L�r>�ty5�c�:��������Pيtc��TT�"(
̖�|�;5�֍��"ƹ�艫�*�ހ�u~|�}zL���7q�g\mgF��ޱ�@�3,R'j��Y`� ��,Gk�-o:oi��m�re������-?�����o�D6�]��tn��/����t��i�b�#,��`��B~�X����4�)J���[�e]��|�f[�4������F�@~�B�ʍB�cV���~�Nw�+B�zwd�!R��0����_�f����/������k#Bd�6�i��#��v��x[Ľ��}����M&��ߢ/&\�!0\�u��
o0s�Ql�� SѴ�26CJ��J-�(�p��wnH�^��[	gg~)ĀN���Q��?o��b�|�v�e��n0����k|E�����o8��י��h�; W-?�kY�]�3���v��|�����N���p/A�%O�0���^�Yi���5T�_�4�W� sY![U�xO����9Ō/�>Ü9@��7Њ9���2`��v� �����E��y�o�7H����?�d���[��`�G��������: ��1xZ�;)I������b8W5�dW����L�#���TE������<iψIg��w�Z�R� ��>?2���!O�o���3��d����+�
�T��� �YX� �k5��Y����eh�%8��e�L��^�8U�[����RΗ඗;�F�,�DK=�K�����SӇu{�(�W=;���;7p�f(��ynk�_��<�����9�+���flHI5��.4�)J�6�4da����u�rww�K��,//�
���]q��U�dQ���Nv�q4c뀱�Э��"��7���w7�S���C��A�f������8���#9̒@�`�mh 魗��-t���E�=�ܜb�7����)���=�'�'��&�_~%t(�����l|4�5�;mm����K��p�E��_eÝs0�:�Ւ��Y�r�䮝�j��������Ty��͗��K�ށ���Sg\i�O��G�s"�E��Xa��Z�e8�u3�n��@G�^�I N����*>��蚷�1Q�FLݝ��%CVs���'&e6����oT���cSb勳� Mg��6y8/�Uf�,���J,K��ݨ�jY�z�%E�Ӟ��;�%A7dv3MfUG�ni*#�
CԚϏڀ�x���b�����	���p��]����m��_�pt�&�j�L'c:9RND�I�L`l;��Ҷ�e���Z%9S8/�?��j��}�Z�H@Yg�*�G�<��?ȗ���b7����-�O.3��JB"b�U�~Sj�����<s�ڸҍ�6]�Rŵ�ɾ{�l�>w_¥��x����P}a�4��WZ�3��TB5$AF��W>�3��l�ݱwi�&~<Z ���EW.'�o;����4��g��d��j�p�����HV"[fff���/�aG�-��ɩ�ʉ�#�Sf�5���O��r-�{���t:T�.]X��R�b���?��΋�nooW���5�̜ P�τ�lT=������~E���*��1�`�ҟP�^7������g�����\�!-�{�o�ӷ�5O��8JZ��e>Zo�Ӫ�ԃ6����te9��B��tj*�B`zr��c�0>��}�ǻ��sL:?8�����u/������d	Ď�z�X�;�������^g>����춾Ɯx�����\5\�)c��7� ��������G�U`�
-��zVR�Oh+).��M�@.L�#�MLLT���*���"@o?@�ܻ�����V�����ϧ2�E��H�I��;��G}D����C�Њ����o�g�y�&�*I�*,rZ�	sI�ύt`�>��Ϟm��[o8YE! �SR	�*�׃��/y� v�2�`[�ƚ��$��(p�7?\�ɾ`���3-֝6y]��Zځ\c�8/������F�zJ��c0�N�,�{�z��2�Q�0�q���Tؓ�G:����Oܜ��k�8�@K����h/��bL�ē�[�me�0��}RJ`���-���sQѹ�Oݺ{*T�t^t5�T|zJRj��ʉ,sb?��T׽_綍(ܛ�j���L�kH���T*;�6S�l���#��[b$ ��I)0��ውR�?9(Kw�
B��T>�L���?�S v���k��I�TlbjF8P�4��v��14�����[v���+��k���8��R����P��_���h4�#i�9���IW�&�N�Ɗ"▛�"�<��HO.M�k�ԉG��I���=,�TD���n�Y�G&~��;񂗳��j�-~s��?���7�'���7��8�Y7P��h�,�K6�%�%��D�C��O`��L!��6��d���V��8����B��8��򪢰�b�i�i�L&N�u�$�a62#�`��N�i���7�G���]� ���؇\&0����_�ϱ�^������������}5kzΙ_g��� ���Wق�}U��f�.܋�p"�w��y��P�~ۦ�g}_g��n�����&�m���~��>L DK3�� m>0!��Gw�%�_sV3��u�P�l�ٟ��ͷ�x�,v�GV:�{"'櫞�T7Z���D���^T�'�Ɨ�V>�,�/��2AD���¬2�{�rPf��e���bn�j���F9Gic!�ɓ��o�ic��,g/KD��E��@�q��� �8ƾ�g�\-�Me��TV(���v�Ut�Cj�c�Q�H��O���'�V�*3#���+��W�:��Y������jX:�[��p}��e����\+L��vL�ǡ���-[c����@A��2؍0@$R{�">AҲ�Z��r�e���"��/b@���`���q3��骹@�e��w��2�����l���.�y2��S������A�,�m��ڗ�S���'e��Axl��C{��kim���~�ʪ帞���3C,v��S ���0��!I����:�����P� ���%1�n�͕D<�-�SZ�"߫f�����GQ[l+p�)|��~O�.���O:��i?�H��fP+���O~���2น�����+��[[#��2��F���'vgpJ�N��"���<|D��Y��(��5W|�6AC���!tSu�5|�+'<�����6H���tϨ������Y��?��:8�d���={e���� ����]H�W曈�! c�J~�mՌ�ԕ]l>�߸�#�	.��]!$��wǂ�"������@�iY��j��c]e�!�<<�u8~��~x�"Z
d�C�,�l��J�6T w��WrҜ �U.W�E�����:�x%E-���z��{��S��G�3�hN|:�g��Tk�:�)�♿w���Z��f	�$�S�N�qhW�v�Ŧ�͡��o��mx�.!Q���������8�
������{���w�Oj��'���T�9�B�����E�:��/�{g�i}�g�/��?m|�	�əŶ�����Gc5��˟7��k��=s��6�.���w�lK���V���C�(H���K~i2�������V�ϯ��zy�'o�jw���<�P�TP"[���u �;8�Z;�::T�G�[~Wyv����9�ف_�p	т�;����W�H��p%�G����Q���EPAZ��o�j�*�B�x��Iw*�z;%X���a���M�b^j ���S�E8��L�d��%ĊD�����sX���k𻀄��1<d�'��=3�A�#�z����j>k��{$)Fh+X3�_Ce��]��AM@z���<B�xKI�Xx�#"Kc��pޠ="���CWr7^f�r�&�\ ��;�z�IX�D�ajn�t��(��E��#z=�����w��Q���KX
���o)n���4˦����ꭻ��y��JV<E4ō���9l�-����TVN����>j�hH���{���A���Q�Ұ�Z�!��Ȑbj\v�ۚD�r�=���.3ŕ>~��Ȇ����+�}���bhc��(�7��Nu����F��yP����%��,��ІDE������D���L���P�U`�6Mc�UW�oZ��̢B/��i3�qX./Mx�Υ�ƶḌ���ڦɝ_T����i���g���$\�_��h|aڧ)�?�g��95��M�8�T����>B�Cj a�;~�)���}�Z��d���Q#�i�FmX�jZ�#@�����츖��R_Pz/�P�T@~�H�Ix�a�?��X$�Kj�Mg���ڵk�:15<a a9a t���w�QՉ�Sjg̏Tn =��֞vmM#�_�����_��`/aLL�\8���Ӄ`��@���9�Ņ����Ye�mO�l*�]x�'oQ��<��-4�ľ��ե���)7@#��/v��⒒z���h<����������k^Y��bM�5=VcE�&�֒o��"��N�`��?���H������m��2C|�n���Ë�\���̳iP��~-/�w9纕��<�f�.��OdP e�=�7���~��KSD[���1×�\c�r��f�;5�Q�V E���w�b�j%/�Q��/?}�O6p��_Ɇ4�gʑM����ƛ��,�ih�^�u���/�T�qP�=�fց�丸����:G~�Ƥ)/�%��e�4TϏKu^!�ѼKW-���<���2m��ψwL�)�������,�����=�V�$�E��΃�m;��Dw53���ܝa�CA��������wj����ȇ���	]QZO �������3#_�N��w��7�a�z]����	�ࠠ��ϟ?����	��)��j���$��U-��AmJ|���m�G��,�p�#kr�����ˁ%ʝ���lA�+$;ʡJ�*�����ǟQ1O�Y��L�؍�5�9^>"�H����0�\t讃miǿ}V��g	!l%-���5-��[@v�������*���g)���,1�(��i�d =�(�{v���DJ,��A��׹���Px�gڨԏ���{�[����h�]�俈��~c�ɩ����="ԟrb�%���QH�����V�z ��c&g���FFF}!@Ӵ�],�w�"�]R�y�L�a�;�p�'�Hq�����Ι��k�����&挱z�S��� n3 0�G�	�0Y��6�DćPb�O˼��N��ߖ��u��	"|����s��O?�	r���<=>~	S
�C� �� �XA��"q�B-�HR��΀��چ���
���}%wOE�ӟ�L�j?�1��[4;��2P�kl�ŀ�HP��G�̙`�DSvPÂ�h�Tא�=�I	Xnj��{y|D�'yflW�8Zs��R�.HA�|�yN+(e6��h*���(��d]c��]j������� �'���S}e5CB��S�� g��eM�w��A�i	cM�_���3wB�5����:D����Y뫕[�KJl/qo_f�[lK��̜�An�|�in�(�Q~�c��f9m������O�+�G�Z	o"c��"�[�tPkY�L�U}f�4	,���:˒�Yb�OXp�<$k���2�;}Q�>@�PjR���}[��~^r��Y~�΃�Nv)��'���~��{���u�3���8�0�h�2�oÚ<2_zؤ�Oi�����SuV޺;��5�;����3��e�+�>�5��3�.:Z�t��%���Dqgg���Ҏ��j9���,~�^ ZDI%�37�|�_��|L ]s��Q}$�}I��U�O�7)�݈��p3�����A�wD$T����`���T*綽gFvF��|�DFKK�Bb툟 �KmA���`�,>+̓�/ׁc-���C��^��w����?M�^���0�Ը!��[P��[����ڹ;�S�yi�I�8��;��� [��CPF�u[��������aP.-S}���4fnz�5��K��]��s�������f���ڐX��u�/Fk�@qBz
�]�`lV�n�m�:�[f(��ù�����\���]0��~^�37"
�@���ן�΀U2�⮫u%@�^ P���'1hEl��o�%�$�6T��YBQ{*�Ea�Y�������{ a���npj�	��넷�/5��)�[�z�$J�}�lQ��L!�}���ߨu��J63ǢZ��g6{�^�i���~'��N�:�]����'���o�U`�{���l�����qcO�>�݀.�e/N}�+�¹B@���6�?J�T7��y�* ��\hY
�Ö~�E�#��1L,������2*� 2�d������@�07Hf-KҜ��Bم��f�T��^�� ��|���i�����l\dkɭ��p�'�Z%@�m"��|�`�?������h@\PAr�@kX'�򧥋��*LrZ��If���8���J��L.���I�S��Y7����#:?�:�ɬ[�4�&/	^9j��S�8�L�`�A<���eI�� T��C��ޔ�����<�}]ϼ�ނ��m+ùw�7��S�X���a�(���b�[a�N���h������i��H��"�� �ςh��
�a��������5�@,Ő��ݥ����Rw#ŏ�1cu�|%��ږ��'|��H>���л`�X������MP��5~ĝ�q���[A�*��	8�6xA:5���������u�����o�:{�K�ڊ�m7�\j�]��!�]%���P2��Kr�M��"�M�vkQ4(M���&]�&+CaL��eH	�眷�����k��s��<���������Ґ��K��M�$��Aw���i{b����`��@-���q$�kq�e!�b���6��4���t�������_�ΗFVg"6S�װ~Ov�hY��?�a/@�|���LFM!$³�#��˿#����332���o� $ j�L�{�!�z��"S3H�T�K_.L�
�vg��;V�Ul�{�\Cgv��!�z$��Xŷ���⮐�v�+V�&�v���u��V�V�N�{r~� �x
hPKR4cC���Ɉz
������Q'�G��J_+4A�\V�e�ҹ��D;w������OY����@jF�~aKw���
�X�R?/T�XH3�5���L$�#�(R�=�.q�?
P�_�&�2�a]Q��(RH�03�~V�{��6����� 矠����I��|�X��Xо��d&/��lc���ެ'LG�%��z�y�����W[�S�rj�{F|�o�W7|��jii�-�;��G�9�@Y^R��yx���Cg�f�#��:O3��kb��H�m�`Ψ����u�1��9���(��npKV�+c`��I�*�\.ٓ'���[����S��D���H��#`:=6?ڕ��d���.6����H�$�4<�m���7�t�,��W-7�����TA�7��i%e���[�6Az�J�V�t|F�	-:��R0�$�(�&S�*�B5p�5��[x� %��|�C�K���z%s�
��0{RZW���Y���k�S��@�y�͠��!�'�%�b���}�m׸���߂k��sZ	�
�~�ȓR���G�TQ�x�/n��,YJ����;�DZ�h}}����:�t�U��ji��_��%xÆ�����hZ�B�mj�]�h�U��r�^䠘��2z��|����Ѫ�����j�d_�n����WK�}�����'a*��E	��9���VVU���}�#(nK��"5�`Ah�U��o���1/�������"�I��}�T��8A�%�ۨ���|e���%��oq6��|l%��+ӆ��ž|�޺�њ'L�F��7���S��[X)GӤ��ܲ;��:���m�L�t?b"l����7MWԉu�0��}���gtRx��ѵ=+Ge���po
Z�D }w5���q����� [:����?��#t�755��:U��->���t���1���dYXm�D����|�� ֢��nk4�@�8��Ldk���N���V��N�����:��H��=NdU
{�A� �Lu�|ŋ��������>�>��Q��.1����;�z�Dښځ��+����+#��y�5��<0߰�H�ڹ�xT���ka�ͧ=�rU-C�1��.���]Ƙ����#��sd� ����<JC)���v��5��c,�f������S�tDai���?dS+��-�'����ԉ�R��r�e�"4*�����G7�� st�o�#4�揦��U�]�wS���(�ܻ� VTGQ�ea��OeБ��?���`�Q��8Zc3�{\��1p�_�U�)�	Y�*���:F��}��)���IB��Y�����ƶ�����@*�Q��W���Z�T�_�xa:���g�)���mu+�%��@�;A�c�͆�;xo���b���c|��96
�(m
la��2ާ���)�@�S�������Ĝ�5-�ãr;�ܟ?8��2����^a@�ru~s��0;���ի��H��L�	�'@����&�FcZ*�詶	].���,Sr�:k�>���s�S�`z';�Wbb":�YA� 2�����ʗ(qgqF�́E�h�N69�ri��P93���[�/��BW�@L:�Zj_�^E��o�X�ʅ���V#�Ɠ�y�+E�A�Z��c��^o�=߰��XA`vbD=��%0�:%�S_���gl�]� \W�ŕ��J]�ڶlҦv���u��C���ZrBT��=w�0����۫]�\H����#,���GO.(1�����C�	iM1�jM���9��9�w_\���a0��Ӗ��Hti�.v4�b������#b�I����>wa�貈��w����[Fi��OO:�wQ(-�����.�*�p[�fϘ�?B�4-�]�-#��a��s^��dGVEch�>�
(���W@�q�L���]!a;x�P捊3Q���x��&sK-�Xl>g>5���p[�ߪ�Ӡ���ʋN���TQַ�0�3\�o^6�Y��YI�#DQQ�#A�ԁ�(3�zmkFq1`,i	 ���%9�F~q[��Őa�����Y �� �y��ǧ�b@Υ�;ܣ������Z�����7�0H��iK�OP�Z�	2Qr�in��~(�w��k���K�09re��f���.9�$d���H��ɱ�'Ն~w�y�V��.H'�Y	�G!�wzݗ?��5���������T��/%W�S��TPi6��'�T'���F��݅���#�	�_Q�ָ�xi��Ps�W��h@�)�{h�whm���zuJ���ܬ�0�]^c��9�o��]?��i�~� %3 ����v�2��I>Ƹgl鷪��g��(VL�Ku�_��Ϯ�M��T�zFa�
Q��hP ����ɗ��g3���mlfڰ��W3�!����c�gT��H���Ooo�x��AȾc���b-��7.H+O.v,���N��㪻h0�ka�Ç�>�����y�FUP���u���В;�!�N�.�
�T:���	����8�u@E��db�¸XWGgj@��N�U����;)e:�u�8��oe�wW,;u���Ө1���
�)��0���7���%�";J��,�,�6���
�x�A&C1�n�I/�0?�mGt�:d�a���V酉���]�[M��Y���y�>�)c����s?��F�+��V49��a���w$V�j�Z���5\�jv�Ü��
i���hٟ��i����<��^�����s���J��]�l����tE���{��)�eG��i����1��`��I��(��Wv���>��Z�v
�HA�Œ�hS��Aȧ���4`e���;_��_Z3S�C�d�Ξ��m������0�.�����#�f(|{M ��T�Z�Q��{�/uȌ��I�!uy)쀬�B�|G^�9�E�r��!�!����N�� =�v��=� k=��f1 ~�*��5ioksKv��GH������|N^ԙ�Ǌ�`X�� Ai�O]d2~t���4$8�%ga��v��i�R	J-�+���q�s���"���u�u2��C��Q~�GC��5J ^�tF�3�W�VF{P
�3.:%�=_p�g�bj�6r�ܬ$�pN��F��B}r�>)��?L�n�Q� ��p|"=�2���E� ��Q6�	ɳ��M��|��o!�*���Ѥk��9���qJ�iK�!����ʼJ�	e�癛��u�$�P<��������
jg�Ƀm�q�hcƨ-�tHS�l�?��5$��\ȱZ����gؼp�"�oԓ�_����(���j-[��°'Q�[h⭡�u���@�҅(�/�̤��$�ѐ�8��j�������Hh�Ը��%��:c�Y��|p]ѳ"4��t�/9�Ȳ�L~U�`l?�§M=ى���=.�nɊ�x�~~S�A�)��	)�L��3���^�i_�ZO��wl����!%�n��=��x��fy쾵K=6�C�J�C���_2�h��p�Tx@.(���G�V�{���9}�m=�!���7vAN��	�"]�4���C/�-��VF-v�]���o���YD����|ބ_P��]��/}�=#���9�:�� Z�h	*�ĕ\�$�Y�zH ��։/8=�H�a#2쾆HV'����u�胶g]���̍�xI�!z��Kڻ�uB�q���h|>��"���<2T����a>-��.�?��=��S��T^�ۇ����]j�w���ť�(�Ԯ�3sD��S�>�x�F�.��h{g��f^r@!\^vgp�'�0U^��și1���j���nI�*�߮�1�к:G�'�3��cB��N\i�`
ŭ=����P��!���pg[ ���N�@�\.��h9DGSn�M,%����D\;�
'&r�/�x���L���^ȕ#��^ˈ�O�kz���\�d�P�_�pT)^[�
Uz��'�D!����Ј����9ROV��ݢ���~��{ٟ��آ*p�xϩ ��c
3�/�4�A*��wAk4�W,=�����<�!��`2J*��!�@�b�
�Ə?/e3�! ��Ͷn3���[WS�<!>�0E�2#�!-XH��~tD�
���mޢ��f��O�v�l��<�d�i#�jM�	e�X�rL�#�X ih-q�;C��6��m9
�S���״T�y�:���βu��%��W�c�����`F"˸���c4z&:vƧ��m/�\������i�Q��o?s�_Q�P���V�9g����eG��/���r���{/揭��w�Y�l�9NM2g��ymǘ�[c#�ё7�oDG�X]�H�"��s�Y�	���T���Dev�q��Ϛ�Ɣ�
2���I H�����X]�`��rp9��?�)[���"u�R������v��R�_�"M K6&|�{]�Q�Ԁ�iP���d3�����
Ъ���G�:ѲL��i���v΀���c\�8@�@�������S흒�-���M��}�h�@�P��Lsǉ��@�Ƨ/�l�M���	�hj�ܹ���:vfW��{A���c���'��T�Q6��*��@x��������=��>Q)jDc9Ʒ�[-���x�c�S\�k]T��>���$.��(Z�q���s4-Ɔ���Y�r���x B�%r��!�S:�?k�
��-0�c�O�&����� ���O����&Hy%.��,:m��J�xCW���x�០}in8ȃ��	��@�$@�՛���[�����:&���;D�?�n��P�� �k{0 �|;Ϭ�q٧�0.0���='��?�w\O~��;�@d��6�Rd���!���lH!�m��9n�Ĕ�%_�qH$2�ᇆ�<�L����m����G�\�(�9m.�Ml<rRMt�˽��{����8�Kjg�4�vB�µ��9��Z��g��w�ƕ-G��)�v�A]WQ<�6R#8B��]=u̓�G@����e=C7�/3� �ė�s����
��9!;�K73sQ�h���f��s���8K�Z��ݻw�8T 7_�6	�ѐAâ���w�!{5��z�	�n��2Ch��.`�0DY�ה����HS�j�-`���8�ܲI ����������xT�J��54,���[���HcI�Sr�A�+_���-�	iXK�ڠ�a?�گͩx�8����m�u�k�g֎���c�w�d�-g�e�w+�	ly������
׼ ��A���A�"IJ��;��>QU��2q��qS���J�u�@�|��D^�F0��f��HuJ����>s���9'Ba~zq�������"�3�b�e;x&!%lk���\��ۏ���YZ'�����7 `��(����w�wG���6�]�#4y����-���_УV�U���p+L��@D�1��d��tWs"���JU�.�l�����h���ϟ:}����-8ܒ:g'�����$ݜ8�興w8S	CW�f�FL�r7z�&����晗OX�sb�o_�ۮRy���� �	�pEEeeT/iMtS�+�q�����c|}�sU��m�����(H�\�[��M�]d�5����b�5�]����+Z.w<�S�M�2�(�*N�1�����h��P'��������M��ȑD��E{
m(�#�o���i^'狎��ks|��h��|hrmC{���o�������I����nx	���ݹ�v%��ճj��{��o���&����3K��x�R��0/��qe:��v�PD��A�|8��{�ft3���lr�щ��!n��J�w)}}}J�nJ��}�R�9��#�@�{p�]n��T��5ϛMB*~�M�|��ZY���u/��߲�_�Z�^sIh��JeC���o� v �pM���5�
�c����z'��~ym�׋�+�@@��/CG�b³U�%b7w0���C���\�)Е�|��&��k�e�*�m-xx�]ځ����3�n����t� �u��K�*����� �}��o� �¾��\Y�yK|	�z+��z����r���=8��j��N m]c����R��V���d���'p�s	2���6��H��9_����Ge%�&1��k����P*T´G ����vn��n�9��;���?@�Z��ܪ���T�Ӯɣ�d�(`9O�J�X��W��9�rǪN=r���Y70�5�+Zx�O/mN[���#��.����8�v��}ϵ)ٷVf�Ǡ�s}�H��f��F��a�@�Id��Ӡ�����G����C���D�U���Є�B�D@!��QX.}�Б�¶Z�m~PK�W���B����d����'�0`��T��w��\"�������&�y#�i2�������c�*�Y8*s�V��㕿�jRl̳$�����D��S�SU�Gk��)�.�ۄJ���`�9����zA��G8��� �G&�$b��9�w#�r�׏ʚI���9zB���:Z��2��~L`�(�D�>�Ԫ��_/K#@^i�"�#��
�&��6��{�	*���H=��I��R�kbЍ�y�)�84򏟻m�⅄�ap꪿�,"�/��M�-��
��O��� �*H���0 J��:�7@�"rr����7�/pOv:�
m`&�&�c�pa�I��mG��x���ԉ�p���
���5_֮��t��9�� I��6��7o>�@p�NM���`�zd<�߶@�T{\Z���XHP�%��u�7�]�9ҟWƝ��Z_�,y�ie�\]�}���m!zPe=�/������m�W�����t�-:a�G^���0{;�5��W��1˂^tޟq_���wlA��{#�F[V�ҹ-N)dGF*Ȩ(L���}^�	�����3���W`bj@+6�^��,�xx�S�x�;��l�:�v�L��@�Z�dǧg�>�T��_�í�tw��?3�GD�*�,p^|\U~^ }��h5���	z�PR����ɳ��d�+�.	3��{��A$�-t)�_;H ��h)����*������ԍ�?G���;hai�0��*O�L��\n�0v��۷�x� ��˹rg�s��/�ޭ��+��A���)����`�t%H�怪�o�oF���G�Ңg�$%%UӨ������U��x�%;�P�}ݱ��'��9�y7�6D�n@U�A��>(��uߤ�/
S�WF2|��?}���l�����Հ�7K72��(��w��Bt�/���8�a�ϴ�W<��Q����n��� ٢�S� z�%�ː*
�������?����6���\r�V5u��A!��� :��PR����G��X)k���tM=�I�$'�c�yИ��]�KB��|�]��5B��m�m��*���5�b�m�|��Æ��+ڍG,h��M���r�O��RY�Zh�M�@��,��G����~'��a�F��Ի������
GB�jEq�#��*-�T��Wo�l�2c)��ro��g��|ǚ����W$�����J��9Bc�E��ָ �X�X�x�Ω����TV�~hM��MN����'�B<�Ğ���I�%��"�d���|A�C{kO@,�T�3PYJ�ڷ'/`0�	�w��M��-�׿#��Pt9i"w|g�����}��H/b�g�i��]E��!��z�W��Ya9�5�{�e�.vqaT��`ٳީ�b��y	�y3���;8�C[�}̩���@�[�vP�]*�)Rf�a���RnM7c�����k`�Gt����e��h�L4�["�z��'��n�; [UlE��q:{AL����>�B彶���Lmk|��ym�ď迊�7���������e�!��=`?1֠�� m��$;��BZ�h�g7�����ĭ�EAe�n���+���
&�y��իj|��(	��b�5��B{�g^�i�n�(���smD�qvno|����KC*�M�gcc�6~�4��I}ڌ���KlP&d�1C��
��;�/����4�-�U�t�t�Kp��:�%��zs�b"�w�`6����_P'}v�w��ڠ=#j(�)N�&�S8�����*�C;���r�پI℣i��'��h��:��.��i��˞�Z�3+����>��==
�R�F��O}���E��ND�*Zڠ}5��-�ͧ@s<�%�U�E&{ OBHѽc|MJ�I�i��m|:=C�<8v^��P2���m�o��n�mv��&�<����,Օ��סʃH�!R���~+F��{�^�Յ�i��
�D2S��N�A�7���xx��;�m^��'��d't�BєqPS��:�3 �s$���1^�j<�Q�	3����E��+�D�bҩ��Ԧ��\;}����M ��'��?���v5U{^�W�`pd��/�ŏ��n4YgŢX�xV��%��h��채2sy��g�>���7�N�S��=�ro_��k��4�v9yO�uvr
������9o�:#3�*IM����9�]�C���C~rwt9�d�'�钠��Y�K7�_f)L~����ۤ���w�Bͮ9Ƕ��Q��	z��c�OU\�yU}{,K��5C�v�������i��ڑW�%;gƮ�H_�q�Gqh5��ؓ��p1'u�C�~�^MLT��!�+?T,o��?v�����5���C�e4�e��=3#?��=��6Xix6/[;g�WH�$R&ZSߏN�D��+^��;�3���u���e�'���`&�m���oB5Qh�D�jr[�����'��W\���&��h��m�5�wzx�c�^��F~MӘqzk�z�9�,~ґg���G�9|_c�[Ԡ��+D+O�D~��[6+�qS��M��FJ��X�؍�C�YrK�#T�UL�
�M�u��΁��hC�Nۈ�����3�@H�������wɜ�,�[���a��M�b<�܀�H��p��o������({�+��B������mbpk}���!��$�GE�2Ԉ�,~��k�E�Sd��W###6x{UQbf~~>��u~1/U#��0 ������r��o2!X
!R�z���	���j��?��C8���*��0s�M]4�;�/�BU�2��ߠ���)e���S�y<���Dj��L�g�Q9�ӟQ��vi�q�*O{W�>�`*r���q�I���u6�Zę*��u��z�ם9/9�4�l�E+�)/<i�{&6����������(g�����-�6� T�5=8j��D ]����{i���f��Gb[�����c��I��	��SOC46�D�i,4*j�Z���^�������Hk��L(��"��ڔ^�	�ƺ;���m�M��������R�q8ףm��N0Ζ����@�L���\�xAV�j��*>�r���/SX	Uo�8�$\��@f�q�oB�t1�K�s":z�J��}�R/K�{�RU6쐈/.iS!�?U��pD�T��XV׻����F�(�R��O�|{�r�����n,i__��jT
_�}�hZ�A�&�Pg3��V�
!x���ՉCFRw����<}��̖\�1�����8�/f���<���)�D.�X�R!2�aɭ-@ޫ�nd�����JT$1t�^�l]�]$�C�
Z�LN`wB;��2;Y�޺� }�P���d��j}$ґs@�{fW��T�N{��S	��� �S_��+i�js�!�M����*��m���޳��dj6$�np�;=,�<���}7�@W9�vĩJ�罄�1�{���7���&x�yԘ�7*꽺�?�4~��W���B��$���7o�,����@��|��[��c�g��~�~CK�v��l�w�j(G�$LWzvr#���)���E��x�MH��n��zC�4���G�iي^ǂd��O��d7�j��"�e���h�f��j�B�m��!�K�U��;#�#a'�j�*�0��ȯ��׳��(I�p��mM����lՂ������0_0�t��PZN�8�a%�_�
r���j�8�7�?緜WKpy���S�"�If���i���S�S�ހx6R*�;<��5U�z��tq������h]�)I��9�Ӱ]8�e�e�M��M��eO�^A��>�:�[=+�d<Zop�p�P������SN��.>�M�������*qA]t{�ɹ�$���:�N@د�`���{K��#ϲ�t�s^�F���%}Gu'{�X@'��c�{dV��'h�cd�&Fٳ�%�I������L��gBKZ�����ai؟�}�+;�?��dz_�Y+�j�[H��M`��\�S�U���vѩ�H�c�)��k�A{��h��S�C��z�Z���hf�T	␭�`u�$�D��ˡ�m�hL����-�����W���[kP^��(�����=�����v{�/Q�����yhM[ܭ2�S�zw�y^x{��vT���ÞR^�TG�3�'}w�a1��>: �N�f��s8S3���NɵlAG�(�f�C���HxZ�2R��ц�����;:H߭�E_9�{X��H���Po�GE.�����#(�"�^���ŶO�z��/��9���u�.�Y��yV0��bj5m�4y�n��&9�����;WT囷�D�7��B1�����s���k�Ӕ�"Ϥ��uʋNU��k� ��1����;3���D<�`:�[�7K������C�E������	��6���W���;j"�1��Jp��
�UT��!4)|��?����_��D��D��ֲ�7�fe>oL�Voϓ����GiJ�=nCv��y��ф���Ԩ��W,=;�������EM
�{s����S� RG�{U�{RU����U�V����I؛��w����N�� '��;�x��3�v-�C6�ɕd>#�s�lL�''`.�]����t���w�q��E���Y���b�m#<��֭R��Y�o�l�q<.�]4�o��w��Cќ�������I Kk�ǃ����qܣDZp����n�ᚭ[�ą��m����n�C_塟�ۑdі.��*��dv�6�r��c�j�rt_�z���W�}�2dꡫ�=Ws�Jp�BWd�Ѥ.��3�ɔ[^ ����h��mnX�K� ����D�
W6��es�:�yz��k]n!�� �q�N�<�0�i��8T�ǘ�'r��@1	q�a������3RhFVS���s��׸��n��=�����2�C�(]����mZ��~�c�A#z�vptt�#*���߇��m4�_�QS&誦� ��-�p*�#�˟��K�kh^i9d���r?B8=*6����$9�յ�z ��&�I����Օ��˱#�<�I��O�k
���rձ��;��Ӟ�)�NY����C����K(����ڠ�Gb�ϑq�U��8|0à=�R�,���=�!�Y�M�XtJ(�h�X���h�^�$ONJϥ�c?�����<��O,�є���`[��?�<��� F�vl�&4E��p�y���Э�-2����%��k�L��"�ſ?�-ɜ�&r�?���M8��M�A�n$���7ԧ�:��z[vS;�\Y����׬^
=P@���,�>��L�X&�_�Z��Tu���W�3��}2Õ="7��]jzX�v�	M�(|o�O,
x>��L���aƔ�H���
�ė�\�;��W9���O�]��Cl�=�5�� ����}l:�+]]]	~� WW�%�3\�AS�"B����݆x4��=�#��0������%}�G4�����C��
���&'������o�OԱ���h���r#�U�@>��h�����(�y��� k�^a� ]�ӟ�~��˰����Q�^!�����0@ލ<��o0v��$���4
f�0���d����fM}��8��n,�)�ŧU���� lt��y�3~�頀7��9i�c?�2����Bȴ�7�H�#eO!��"��"IZѠ�2�_�&W���7o���3��x&4���Hcdu���� ��G�߿OV:u��!R�!�bChd�Oi��|��	lL�#?�XuMP�O؂��|>o���=�s~�%x�+'u)�:�$l�o4{xxT�`����{����24�w8���|�K�2�G?;��	8���nN�������^�|AHӿ|���l"jz�K��"��W��@����O�ɜ"����Y{m9�3J��&9~x�"SD�h���1~1��2��4�����U_H=�$��/���/��3j*�3��*7��4�J�.�|/��K��.��7<���z���~RuU����K�v0ޢbִ'i9�rf��g�.����A������m�8�=�(�!y�!���hᎼ��=fs@�*;��.�U��fS��~y(&�<N�I�ܴՓ8�>�f�Rb�%hn!n�A4�wE�&z lEcĸ��w���@��H��`a��W�n��0�C�$	��5�~��C�'�ji�}�v�xIa
)�'ZvgDՁ�&w��B����æv�x ʝ�٢�c��6�O8vN�b�0��A>���|��3�",��mE+�UO}{�J��Ҥ(���{<��@9rR��L)Z��q�L�H\�����*l�_`�V̵K�+m�f�e���h����ÌM��J�GR�w}��\ׁ4��1��W��C1D�pV>���p��=��:���T��(N�5"�D�}��Xxl3�4��ox��j'{��?��ag�����sT�����n7{����k�M0-J9*���l^Z��_��}�˗�'o�%J�Ю(��cSI���
��6�h� ]��{ܗ�&�~|���:��;ft�9Ry���/�5J�E������VM|�$v���S��@1f'BW���T�k�G��͞���K�P�� �Z$B����ۣ^	��uD�sKT��}����t��DS\��t��8�2�W�&�2&|����9�|�:{�Z\O�LLJ�1G�Q�s�\���G��'�j!n�(Q�,�$�<#�y��E�B�RW�DH���>.;L� �p0+x���\-D¹Â���9��b���6u-�#l�Q;q�����G㶚�Ł`�'2jԶ��
��,H�T�9��/\r�dEL~U,�R��Aѡ�7��%r8��u��D�&�-���ы��#� ��t�3�d�%��{��a�Uh�(��8A.7i��v�)xޫ�7@бԈP�lo����8h)E�%�mW�g�+;��th�x�]-J���Uj9{T����P�q����/t����t3����&vj]7y+_�=0�R�s~	h ?�؛܀KQ���G�Ll��|������/�.�{I�@�ܳy��uاȀ؀�6��}�ҵ�����
H�(n���{�����ע&��j\�j����$�~��|}�=�rp!��@OS�p�@���2̅:�e%���%��B�������nD�k�,=]@���}�i=L��-���� �;�����wH�����Fo�t�736�ʱ/��MLG�.�=��r���s�(�߼qꔑWK�l_�f4cn�#�e���k�����h�ɗ�t�w�5%xFxM����j�����&Z!��AX�tA�`˛�1q���^�X9�/��i��U���Ǎi���3�/$�6Z&�<#+k�Ͳ�ծ���=:�6���+h����;>�v�L�!�S����Κ�(wlr�z����E�G���{�ծ�y+;0A���g��><��&	�(���H/��J�F�$#Q�&cպ�Ca���1�:�2}���>��V��o�n�=u��O�6} ���>>>3�����f�,�`���"�B;�;~^�J��M$-~�~w���=�����9��\����Y�}!����8s�%�h����q}����(�6XM�mMie%�n{����r�M�щX^a�(�6L�n0�/}D�!�)���8e�Gn��#	�l�{\%Ϗ�� s}�j?�m$U�t��c�ܩ_ �^�L��y(�p}l���nz�R�iU����HK��ڋ�C9Ż�0��E�q���Τ�%�h}~���Y�:0֊���X5l.F�G� �s���=1	����91�L������44��D{��'T����Z��^���`<JQ�+a�!��Ρ#�L�`���d�]$��&G�<%	��FMM���Ĩ���l D�75���nBkt�:B��'����0�>�;ohhz�'x��d鯩=F�����]g�K5�x�^�ul�ϣi�9�*Љ���W�Z�ć7���nu(fب����W��X�l�����P���}g��.y�\�Җ�C��zn�T��ccc����2�|T;4���C_��'CB�νV��3T*������|�����=f������jK��B��hZ�n�ki�.�ѡ�mgFބ��T���LӦ��)��_��s��r�n�ЀΡ��C멝zy�=��Ao�����lg��N]F�g������R[�[�:�?-/<��{`��i9�R1��A�<������0I���V\�:i�R��T�"F����g�'x��6�g��o������ڗs3#^{  p��+/�h�8>�h��a֞Pb�.Ȫ3Ҟ�X�q��-~�"{;x�L����[F��kuN�^��Z�M8�fה�OB&�������t��z�:_r���_�����3���S����
Y��;M:EK)����S�Mm�^;�~[���.�nE�0T��0��mO���ݘ�b��.��/�%䦣2���w0b��������?�o��H�K�jy%K�Τ�k�'ԳF��`D`��g"��B)3��ee�34����jMiv��W7����h�(�PZN,�ptd2)�(�+�nv���X����=Z�߱v�
pf&8�qP��o#F��$6�Y]�Z��}��}��I[��+��xn)��hC��9e��kߧ��U�0�t_;��f���h9x\�k\��|Q�>}�Pp�f<rF���.BQP�J�\��d���Ka�]-J% ��T��2يk@�\�,2��Q�_������A1��g��D)�*�yC��/�	i�wV�$��4g��p���ݟր뉶 �𧦕ձ�U;!HR�]L	Y���}m������3-�����wO<��n�i��jW՚����}�
���$kDQ��^�J�<J����K[ƣ��z�u2!�w�q*f��߇��KZ��Q�P�	�ড়P1� OF�L�u�NL�}�����Ʋ�5��Q*�~�dz^�f�q�{F�<�3�[����B ��r�C#r5�o�^	�g����!�dx��-��PL݅�>}4�x z|��M~�X�$Z��� D���b3xHZ<^���ŜߝX�LvP0�ۢ�у����|��v�s] >-�P�Nk�5g�­kK�����~�#}X��q�ͮ��>��[�%g3�4=������{���5Ԙ.���
��������Z�:�,�O@��q�'��ح�y��I�:Ѓ�z�.2�l6�����I��[d�-��&� ��j��Z]1��Sy�p�ƕ�;a�[�q�ѤL������<�5��~ק�GM�8mn���_�l&��-����_H /�����L�����k�)ʘ�߫���z�SyWHT���q�C��X&q�}��uk��J��ϕ�~K�A�PL-��lWd^ý]on��8�T.��~d���1�(�(d�S�&Ɋz��c/��W�<틈aQס7� �-F��m	$�͗R��$>���Ӓz�^��K�xe��W�W9��_S��Y�`��3��|���㹖ȖD�� Gt���QV�: ���R�P���=��:��)
}�<����ѡ�o�_k'&&lJ����i<k=�n%�D�6��l�Y5����+���s�BA2:��z��W���Y���*.�utC_f�?��
�~�)��P%�K���pV����=��"'�EVw�x�v��}j� �Gvy�t�o[c���,���Tn�⢀&U��Z]Q�rސBV��W�,���)ˀ!�c��2���01��'�($�I^�����R)A��@*\َ{CE����7 �+�{�7ܕ�(+~>�jG�υ�'<Xum�f+PE�-���^�΄쟸A�p��3Q/��}�������S^��Ρ���ה��k�Z��0�Ïo�Ү��s
_�����*B��Z�4���3�,.Љ�,��%��o���������sI�̔Bg�*̤��yڷ��U��� >�*Z\a\3k�?����V硿�oE�������M8���K�^��#�¥�]��v�`�:���m��Ya��휣�b�R^�i]wD���Y(-1��h"d�{m����5k�U�������Hw"'��7�`<��z������D�O������~>.����#�ﴞ�_�'�����!���F`۬�]1*�)(WIY-+B��2�rL/� ��c>�N�`��&��e\b!	�����ߥ�6�(�l\�v�tq��/���5���xe�*j��)�����p�^���Hs@L-ߐd��C�����
k�'m��]�[Y�^0VO�e@ *]~ ��5���"�	���)��j���Z-Pve$r��"c��Q��v����ޑg���)c~���p��|z�H��Y>|V�K>>nG�v�t�P��Q�T^�2�۶����
�1�/T C���f,��b�� Ib�Cq�Q�7��^�,�K��Z����if� 竳�FqX��S�*Z�,����c����҆<xSO�p>,grz���w?(܀H�
e�����[��|�["${����!r�Άƀv�be�W �-���������3gu$��/�j1`u��q��?����bE2�P� �f���Id��B):��N ����+�}�
k�6��f����v5>�靁H��@˫�9�P	���(�XB�Z!���[�jXJ<�]��`�Ѡ)�v���l,F��I�)��| ��@W�1j>c~���ys'��i��'�M6�9����?!0�C$�8E���D�(��a]X ;p���"�3�__m��`��3.]zO��£iJ#�^�C����΋��=�[���AyX��?+Zě��74��*���4�:�[G%�s�y���M��|��(�m�j�� aԞ=�4�0���r;�3��<��X�`TZ������L��m��@�{5Z^���Rؗ)�ԏ�l�ދgO�O�t��lE�y=��U2;y)�4���^5.^�%��,�G'&� �ٯ�Y8�s���/{�E(lp, �������F�뽇{
ʱ�s�㹅{�+�S�ˆ$��B(0����]�����|wr��,��~�v�=�'A���y�,���}����0�n�|�u��+�D�u���çQ*g!�Af?"}���)E8!$�W#����e;�T<ic���>�O+�N�uEX��F@��\�Z�E�4�ߌp���!��ЏӦ����9AO����(����8����/ �&������Kjg~�(�Mgo��R&�WҰ^��^m���S`�:�f�{|:ς@�-�{�.�D`�?�� �mF�������aB	z����Y1[��lG%�r�D��Z��0�@��:�[���[���M���:B��\n�7�l�N�i�}4���3�H��!��������߀�tm/�k|��Њv3䡜>/x���|U��A!f#��ku]��jas�F���������0Y�9�xZӁ���-�q_Ѫݑ��適>�ղ���l�#����O᎟d=��O=����i����y��B�>�ĪO��?�������<Uσ;�T	ݻ�+fg����mL4�@4��I���L� �3�d���
���2�#g���?a�Ⱦ_e�9���V�54��Q;yG��/j"�H�ajg+�՗�@�C�k�V�nuZ�f���_0����f7��4S�E��$�1q��e,��#�1�r�n�S]VV������I��`��O�Eu�:j�%�F.<�C}x�Զ���	s�r�5�oA����Q\�%��6Bh���wA-��l��� �8!�g$	�&��d�����X+�+����>S�xd@���\E~�Q������̡�#9R��}��������}�F?�NϞ	_�6�|EtȻG����[*fȸ�Z��J�l�+1�:-	��u��0�gB�hFT�@���kh��1{��Ay�7�(�'��Jz�������ձvLL�`�xTr�#}��|oMħ�zy�3Hu�O[�@SH=n��rq�E��m���Z^�2L�O��i8���zm��~M��Ѧk�D�/\��"���ˊ�A\��'��:��P�l
s�� '�^�n@�\9�>y�=p�+c�����r�cͼ���>b�Cp�mA�?���W��B"�J���>�5�p	����ȿR||��_��5�]�Fs��hÉ���A�!�RY�l����N���7	Mm2.������|��0K^��Ð`>�1.� �.�~�a�Zi�-��2���x{mJn�*�束�O��H_l� ���'A���E�v0���3W@�נ�׃!<t.�垺{b��ub.�W����ne��&�A��K	�9ϐi�$_U�C��c�� |2�\���Q�H�0�g�ΚC�J i5�DW���#�q�xᳲ�� ���zv=>Nh��c��ߕ�����j�4?�������-i-�I����d.�����Tc�dVa�w1~�=�9�:8��1=vM�l���(��x��1kroHA��p�#��mt��F�g���U�w	Ew�Yn�U�!����>j'h��r='롸N��mvlI�����k���:���Qu�å����d���{޶I����s��'�����S{����F?瞅���S�(=�bTV��.]A=I��n����YzV����|���2n�:�ѼQ�Y�&�#{UR*H�S�q������U<���-��@��-{ݬ"���v>y��fX(np��<���W�N�ko�CWK+-�E7F�H�ӂP�����+�[X1Ÿ��kd%�����SΨ��d�#WO~(��EΝ�?Z�oٌp�t�T#8�`3{�0�J�����d`Hq![=�<��r�!�+��W]�)eS-��;z�<��,TҼ,~���Ktg ��ڳ�o�+��J�Y]]��`�v?��*@��pU����ޟ�S�����4h$�Q�J%
E�ШdHi3��%)�$TN���쎐�:Bbۆb2O��Y�Y�:�߿���^�w��~����p߯�u��{����%��K�o��}ς���PͅKKP߇�b�XC�Jh,�J��a'M�S)��k7���J:�|�f&�O[��h����
�Do`E�%�Ⱥr"���y�u�ڮ�i�L���řV\K��H�E�dIC��4�1ִrW�Ps����9aM����{%�Y�]D��ޕMu�jY�[q�Խ ��]�;�m)�F��!�/�
��j#q#ٺ���Q��y�vXta��)���f]&#���É`�8�M__!�.ӌlxB�'o���\�ՖEtdІ5��N��ʝ�'���=�],v�tw���Hl�K*��t�ZD9���t�0�#(ԓ���ͦ�1��H�:� T��t���:���,OgJ�h�#�1��V%ئ�
�]+H!3/�������Gtb�:$t����ŘH�6���gf�4A��٦s�m`���R��:Y�]�ҧ_9gpVk���\-q�?�81����������#���w�%�C8�FS�PA�2Q�ѓ����R�k����&Ժ�LS�B����v��#؃͋�A$���1Ã�:��9_��^�g��k��<?_��I�Θ9x i�.�Y���+�9@g��Ϡ�x�(��3��$�&�v$>y@�I�!�e�fG�ڮV�%��IlN����W��O�C�Ğ'���?`h�Ǔ��z}+v�=�]��i��Zsf����[E�_�����b����3��
�Z�x�X�y��a�-Oi��jc�f�}m�tU�0�2���)��T�X�`1�v�s@Q�(:���XD|��@g/��y�j��"ZF0����/��C����G%��_�?dr~�$v�r1ֺ�a����&@�����`YR��ŏ��%��ʣ�=�6 2 zBm-NΆa#���H�e��,B]���W�g���I
'���.��'�b�Dg�k��e�/(*���ق�����8�Qq�V��ںM��)�,η����\v�����ӳS�.�������'d�X��+DP?ڸ<�jw^�,��S�>�A��c���i4�%�y�F��#��3a��	8�)lSU`m�3.(�,S1X�4���U[}���.�7y�>�̾�_���5��:��j���4dp ���Do5�[d�2F�c�"1�Vq�j�cdb�ٸ��
J�E¿�z���3�׍�3�z�1i0��]p�U2��q��H~S�B�B�w�G�"�
��*�{�?f��h#�������	���m8t
������M��0,xj^�<�e�#Rǯ��R*�qV��4B���]�[��l�:x�ʻ�Y�Q��y{�L�2�}��X�u�v�	���}'P�������@I=ϿɈL���O���Y
�(�<����M��C[�T�z�Lߊ���`��H�����DL�#�FFze�H�
�2���@Q�7���B�Io��!J�X��b��Iڴ��ӹ�Q/iS>Q�_�0��=Bh��i(�Pi��T+��#�i��~~~��*_����cۨ�w� �)9?�G��e(O���Rw�&:���=!���=qd<,�zx�2e�xł�2'O(�^�!׊��Ǔ楞��:� V������j���E��O�Ǒ��H��]�&�T���V������)���X�Q9J��-���ߝ���h'E��Wgo�J%� Ü�����y����%����8#�$��viT����y+!����rG��VA��I�E$��n��n�.�S;�&����Y*�x������ۙ��'���kb']��-t�J�
��~�%���7�˝�;��o4���Ź2՟�W��ؗ�L�����XG�|Mw�^w6oq(wP�K����(h�/_vOs������f����ʇOt<�y��l��t���ӵ�S�/+2ӧp��7+�/w1�z�/lMc�����}Ip���'� Ǫ�wH�5���>J|�蓶���5�Yo��㐡��t3�\��ʽRMK.�ǂ	e�m^�_}�7!�Us!Π�o�ܹ�f�f�P�:�f!����cT=P>��u([C:e����o:�2��;`U,�υ�+�^�ki�2��2���A���]�m�Apr;��>gǊ��+���ΰa؆��7������m�uO��������_HP��c��>�v��R`�o��l�C�����cLdz3Ф6r�8՝��-|.)����KX!ո0]����E�7N��-��=ޝ���P-�Kq�<����;+,�$b����ҁ�錓HE+ksH�������w��fd��$��˕'�?�ܫC�|S,���CNx�y���N�Ng)9��K�Kc���o�瀧���.�?�3լ��'��u����+����JNE�#A�x?##C����=�(�ؗ���w�~S��E�t�K}}=i.�?����c��1�� �GCV�e���_�������@��=E�(�m��/��h
�.�R�JZ6�	9̆�iCgg�OۂC+�B|}ۖ3����V�����X���1t�be�h���R���	%�ju��� ^t����`���ӵ^������9�.�Q����Yfn�&j�݇T��j�H{V���TL,�Q-M=�!s5�C-�����ɔ��<B�c�I�)�g'g$��1���o���k��	J]��<�l(9���C����6\���	�-l�z���>^��9�ӊM�/��%�=��lxD:����ṛ���կ,W�k�P�]�~���ٽ�=n�ߪ8��j���˛�w���\!U���Ef���2̚v�yυV1�[f�drQ����yv��u���̯��?w%�)��+�;����]���]���j�ΣL��Xyl���������i��xC0�\�]�]��&(��F>���x;0����qΏ��狘Umtx��`|�����Vg�@�B��y�)��ܼ�,�L���W�hP�Ӓ�?����s�Sا�� Ã���\�˝oFz�)(W�ǐ�-%�ۮ.'�}ؒ��_lE�$��=��|Y��*��oM�o/�`��+M��\'�'�w�W�@>�qt����ѽ�Qظ]N��a�=[�6���xԼ���>����P�X�0�5曆����v�w%1ӵ�{|�m�h+��o5!�_K��P)Ͱ�9��9�n� ���WY���pִ������YC���R���%ў����o6gM�L!����T�Pp[�����o������k�G#� l��:�j����n'�C����2���� �ڌ������8'f�L�Ȝ�f�r������{<F�r}�L��7�4���x�����9!��� #���BE(�ր�����辅��~ju@�%`�j�풙d|m���d�lS>���#s�m�fΥo���M93\�'ݍ���n�Si�֮/�%�&џ����Hִ����!oB�y���Q�zJxq5DvcP۴C��9ūq��7�t�>J�_����(����8H�ڸ�S�>y��H���������t�b��bF5Ѷf�R{�4v�_�K+��P|$Z�m�;ў>�f�]_8����X�f�1�IK�y2��}�>��*]�«��-�	W��:-`�M�Hv��F!��HS�&b�8%&Q�̪��[�pS�v�o6�l�\��ʜ�v����N�������C���BA��Y��#v��SY��⼇>�}pZqY�Q8�8��j��BKc)S�A��@��^�����]0�O��s��;���]�QNv�ei��)ĈY��ZϚan�꧓|�.՗�J�:wLĲ��	ɢ�?�q
z�"�[0��]��1g¢r�k�/0P ���4�fF��M���I:��WGQ�Yf�{ �mC�𯴡&A�CXE����GCv�.,&R4�<�1e�tљ��e�2������u>FN�	��WG/�a��򇶢����>^�>��y����`M�TmqP̊�n�W�q������?�1��;��v�	,L�~d�.sJ��(E ����5u�EQ�fY���i��:�`}\��T4C�c#���v��w����Œ�J�p�!(�q�c���Y!����Lm��e� "��$I$UXm�d���&$�@	�K�����c�<j��W�>��̌%�5�J��	 ���ӟ"e7��ƒ�;qХ4YԱ�㥯�P�@ˊ��)&�ksϱA�A�r�K��"�������@b��>F �O�����~3�)��9�`���ǗL�9��y�{�A2ω����~> ���k��m�
ʘ �m���BL��;�.šXsoddĂ@w �b����?�:=�ZeV|{�)���]K[.!��_���"܉}S	�B��`��*�G�X6�h%�����G(dv�y��N����9���u2�ξ)���=�6'�_P�	B39�׆��1����<�R����g���'�pS�
�;S^���[�+w���K'm}7��"&l�Ӽ��A�R�N� �v�X;u�l��֧(�#{�^,��5;�Q4��l�-$��x�sw��������]�>^�y����,��$�(O��9�ƿ��=F�K��Y%Sf�C3������$��e�{�W{8��im�}�p	���V/|�KK�ɓi��]qj�L�5���.#�5���|$%&s�=��C�1� ����Z~%�2O��+��$c�Z��i����s;�*�,�	B��rR[������KBii6۸4��8��)It[�(�4�F�;��&�5b�kh#M�3��(���wn�>lZW��?:D,X`�"�H#z:�|\���{S5�Ub����b;�����\]I5͝�װqF;e
�8Zg���X_�@��6;��HEWC�<2�(:������~�ߙ�KO�����yyy��"47�$���������0��[��[��Ry�h���F��
E��;�f�>����@�x�2���S�^�XJ '��`!�d�Sʚ�� ��ϋ6<��uo��)��J����u����6�K�o��-��%�����K>�$��}.�����o��-��%�߿d]Χ��d��8�k�,شtQ�k	�w��'?�9���NP����l��b��/�G���8�E�b��դO]���YS����I3�a������N��l��_��=w�=����_�����Ԅ��<�x�΢G�9�X�x���xYeŻ�p���lʷ��Lr�W���'��+�cC3Uߥu3� ��X��%⋞k�r0m���F����+�
�/o�Qx���H����=�0����Ig��I��Օ(D���u�'����3̓��ȋ�&o��}7uss�����L�n�1���ϒxmК�N�:l��������L�M��͇$Ѓm��.%��1~�;��Ï�S�u/�X9�<��kj'���5�r-�G�q�o�+**X��sx'N\O�u���fr�����|�����!�x���߾~}��X;���e����	�h�Փ��O<w�ɝ���>������!��XK���&�`����yy'���S�=_
�ք�������'��3�6�T�VR���/�?WH}nP���G�w�
�M�7|`ZC���hu����)\+#q��;�sVV[�f�]mt�'�����c��]�����KľL�q����޾w���n5��8�u���())��}l���>�����<��%�t&O���Ŗ��$��Dٽ+��s�c
��z۸F�]+�g	�0�����ݓ5�L�z2w��Sh�ME�*�՗s'����Z���m>��K�~���4U%��d�](E'�<����Ν����Y@��e�zI�K&����`�/x��X%��ܖxhZ�&/#����G���@�}_G�����/gg�E��1�8�v聘�ĜOn�x5U��[kIݲسg���7K���{�ʪ�P�j �h���ۄx��U�yRNJ��|֫�3rK˼���HI��K��+6OP
*��W���}IYY�>�٢;M�:�}�$��1�U��F@�͍����1#���l{�
�]���RZ �=�j�٪��u��a�����x����.��'$$�$���i3�6��"�����ay�w�=�<�#��t��|����P��P��5�p���YƑ/⍿��P�T��L"W��^�H�h��}�����¢d�]�=��t�Ѹr��"u-��K�
���N�
�	�]�FX����z�t:f�0�3yx�Ҽ��ɵ�����������W
��S2k\�򭶬�Mc�QV��t�o�uN�Hԇ�"��5	��ș qCR�����Ż�Yj�l�c֬Ys+�Ħ��� �`9�$�G^�g�2�Y�y}ʑ�	,� Iu8��j�+ٙ�����;�(��}��á�D���,z�֚彽�1�!����ew�0?|�p���=d��5�j�[Z���;1P�rQQ����_��"�R��h>�'�ؓ����g��QZVV������� Y�,�Nۯ��C�����E��x4�^�xx�9Ȅ�܉����x����v)H�7 O���d_y A�	5gq]��V�%T�-n�U v8�i��ݻw
�`�����H?	���e�4������ڊ�F�U�gj;;;���y������,�r�'D�ꙃ	N*�$I�l�䜳�@���TwVXX��E�~g �/�P�=f���C�s��ȓ�ʩ������ɰ��k��ҹ�o5����K��8�@���Y��\>����v�)l.�6ـ� ��l$"a�H�����>8!^�q�"�2���ֹ����꠨�"��و0���6�����[�D��kп�������UZ0e�jEp��Pҫ�4�*�77���;�(�����_o������&3D ���_�x�K��no�N����>H�J���)������V[FH:u�C����g�G^nt�����_�ǲ@Ą(��9�HBy���c�Zw�\i���颦I�y�!)���l�o�o)�eOw O��׸�e�p]�V�U'F�}����`u�h��j#h�8aE��\��I��
9A����~�@4�u��ȠT�AX<�a�?}}}e���5i(�ӭD
�Ҋ�XND��F��g�\q�;��?u�#Ȟ_ӧT�^��F�D�/O,vPШIZ�0$��XG:B��s���ψ���G�������\�Ȭ���Z�S8Jڎ�6
OĔ��p�3���3簦�8�����`_�l�$�����K=��K��Y����zezhl��� ^DP糳�S��?��z|>��
�����+㇓kX��<�Y@���T��c�����	3�F�ӹ�\�����dw?͇��SrEݜ�?)������X��X�|#��8 .H��.z���ϟ>�vR�%t�p�51�c�%�������s0���'���NЯ���Ќ	�Z����_�F[
O�6�a����0o����(i@n��H��Z�o	z9-6+s�/4S�U���l&(9���!�-_JN<���%H�6��
��Z��Ʒ�ՈWx08��Z�=�����	�����ju0����~��[|IFٖ��������|�>b����?%�>e	.�qV���>��V��Rɾ��Pv��̿�P�$� ��{&P<�d2&R��ƙ�!�(h�M7>"�=l��F�;�NG�1�"#�4+O������=_A��Z��KI��F��0z�\r)��V�t�^<ovtt|x�j��ϗ�9c/�:�Iݸ0�&-H\��SI<����j��ӳ�=]]\��IjD߲�]_�(��-�l�PeY�_����3�a-Mf��|(`��� ��<�{b��5
�q�[�)�9���<��]X$��HpǕ��ֺy�~!sI@A���_�&h_bz>D"C\C�za�����P�BfZF��cFF�6�#��8~i%?��}~����BHpH\k���˗焊'B "<�㡥�l2����u=z.��W����B0"W^k�����߲�ju=BGuʈ�|�߬A< �?P<�3���2]P�z+[�����U�m;���o�&:V�	e]�_[	�J���u�\,�E[ֳ2��4S�ѭ�����͑���D�e�SI^y�
Ƒ�e>h%��ڬ�0J�c�Z�٫x���0�[Éߕ�:q8�7��
�: ����ε3@?6-�hu��"�����X��y�p|����=�`��f�sX _�G���sQܐ�3ӎ\��O���5�m�v�@1�����7h��a'lE��`����Y4=h�C���	�$��P���Ȁ�%LTM"{��v�#��R��i�lBO���S���nd����c��pҘ�U��ЎL�M%g�h���� Z��v s~�\ �K�Q�O@ �m����J��@�/�<�qߴ�w�\n�Q�AS���|�o� �@����3}�RG@蜟�t �PCÉR%�A���N��p��Zm����D~P��x��6�0�X����$L����P߉��kyAb��SS����$$?w���E��-m�D ����ƴ8�Լ6�p/mQ9�b;��S� ­�ʪ�<��%��,eS�<���+��\4�301�<���f�!F�Ӏ��|��K;ہ��������G�Y�ś+a̡���'��$�SVvp8�l�� ��fNc?+##Î�7tP�1�pI�M����8��|X�q7��p�f8s��������1ϒ��o ��^^^Q � (ـ�,(���\%��m8z{��K�){{{;gg����b�yN�x��#vt,��U�|�! �K'�}�&�P'Z�PE1p�t*����u-GLjz����ȴz�'���T~��~���Qd ���|T��\N�-�̾Π%>�.k�d���5B�p%�A�b���<Fm�LiZ���\���5'�[�Ò�eAAA{F}x�S��C2�(-�$K�s����x��1	�7������gTy��
�4��F|��Y#��8`�����	�Y �g���sEX�j ����X��USR�K��Z�3��@q�z}P?ꛠ
e����e��_5�����j���L>�&�/P���[s�.�1捞6�w����ETDd"b��H�p[#
��䱱����p[,�@heq��+9g�8�UI�;Q��`pĆ�y���hsf����nNN���C�M��p�7>^�� �Ċ[Ʈ +;���L`Ts��MM�
�\�)��>yG�T�t�)�g�p��_��^K�t޸��y�>�tC�'x���֞#)%�IƝ����?Y9d����@��m��x�u8��V���Y��f6���ڞ�\"XsJ����%XM�f�!BΌ����?`l�Wu���(k5Z���'p�ף�f�&��!dw��[WX�BLG>�_r3���-?:D��!=�PE�e��w��������=���}۷����"�1�_~ �DSq&Y���:VHܴ�8��&t�F�y��g�-~d�%>��ضe��%��P�YXX����1=��?z
�)` ����BjY�tYY���hޣ�,�f�'�I,C� EFH�tΨ]FR�,/�b�D����͓��������3O�bWW/�
N}I�Kh�@q^b�&b)S������\mVP���Q��C���R��,/����]ڰ�����d��k��Czu��@PN2��8<KQ{�k:�O���0gB����|*\�/9��28��1n��MT�G�L�^� QU:�WUH�d@M>m���"͎���/��ֲ�xВ�ɏ8�GQd��gl�l�M���6O�t$7(B$)�?�VX<��_�I*q�'O�o.	+��&�Eo���q���#VA]Э{� 1=*��7���tz[��W-/y�% 吺H��#\�'Z=�<}]�f/R�)ݍᤴ]�.�1MnO%�8�+���9V�a}Z.6�k�__�H8��gh��Юh�#�:(�Qp�[�,��V�At[ �������}�
Tx%���豦��ka ���"V�5�^�SO0�J���9IV(��r���Ff;�<��K6:�&ЋU_�F���t>J
 wW��w�R��y3Pdځ�h5R�ǝqrrzO�l�4b�jM��.��[g�*"�"E�T�֊@��X�j9�N�q��2��Zq�j�	!wb
�c� m������<��K���p[&��j�� �yJ�r_���	����a�c\�P���#w�(#��8!iZ-��8���G���5>�Yپ_t��ĸ��xv�����Pe���Z��ə2�Q&�����[�?����{x�}�4�b��A+��C=h�C��`w(½���c�PW�����eQ���i��k�3�S�1���SS?Q�v�0!��oUD�2��yyy�'��o aXS��܃�e���4���Y�A�o�6���6���Ci'���;�##�j&�BB�c�;::��������^�)�-�ide�_ī�q�����6@��$K (�Q9߿U%eDEE����S'���M����42[���@���W.�����>2`ooo8�D��Z�/Xs�eJu~G�q]'䖖��s���x^~~~&��<����VWWǐ���(��	�[W�e���ͳ��/����8J=ej�/�A Pt%U����a��x�����J��$:��vǓ4�+��(a���S�œy�'z�	&9��� `�#ěڈg�!�Y���8	�!!!7�S@3��pg��	��ё`"@�&�~y��w��PHyrJ6���r��ǜ��B�ĨD�)){(<�6L��R����M-�Pϲ:�:,���b��U/�rw����ꉊ��Kӣ��'�j�~%"<(Z@:#�<L�.��#e�l�"n���h�9��[`,�Yl�ᘱ+C�w�v��c�qU�ZS/�a�I�s�.��?�k�iϞ��h��p�S��p�r�3��3��3><��F7Q���y�����.���!ƭ��_� �>�$w(C�B:�viA��Lv��rd)��������B��&����Ԡ�FQ���Tdd$���@�����X,���*a(�R$_���ܰ*y��4t��	����H>�r�Jf���mkKX^LLL���F��Jj��� ����	a�e8q�L�np�]g�?��`��.�o�}||0�1S�Sj=�t��8*! 	͉ll8�p]��L���|�O�ƃ�\��"������)D�IS�V��Q�>�ycw*΢���l+
��޽k���1#��J&Ҥd�1�'Nl��	B=����b�<�?�`u26>�Y�m�܅�x�:���<�	>�|�\龸p�_.��}vt��_�����/�Y�����}i���+^|8�W���T��{�$2<<gC��8�t�НOt�@�V8d�>�����[�Ŕ��^���?��p�9U
�[ww�a<���ד�Iii��N�H�w�*+QJQ��fy�'T&����f�l��f�A�6KrÆ���ʄh�Ș]L���29���"��f[AE��왭H�����$�u�)�2 6�>��{	6���%ǌ���-��(,$)�P3���144D�*�P��l�'�рqU���fnnNOy�2]K�!(����^�����e�C���'FRa%͖�2��Z��g��@{a`��šq��]���ߠ.Ȓ�T�݋'��ت�����o��}J�N�X�c`$�ܥ���
tk�H@������X�q��o$ZgS7���[F}P�Ћ�n�@�l����
�4�y:�]I	�ܓ���ʪ�	dޥ=�!�yU��u6��POS�hUU��E�%��~w�����v��b��u��l�0)��������Ap�^j[�/x^��<�Adt�X����y�v�eFHH�+����i�e�}� �Y�ٍ���;���*����("� � �
<���@!�.E8ST
g(����h����^YY��`0DvGiwrJ��|<*�s�ܘ���`��*咖���Rge�m���xg-�e=?�^*VR�p-c��ى�X��,���A	��0���̰���qn7J�S(�~Qeq�H ��@L�0����[�B��kEd��������* �����MފA���a8���;
�vy�`�VBBB�Zu�����zks�y
b��
��;)�q]�T���ɭ��t4�P���0�ɭK�:
[��$G���rѓ�[����B
=���(_���s�b��R���&3�(r_��h�A��o�⢿����Le
P&���5VVVw�\�}�H�c~/��u(�|VXX�	�&���@ſr�d��&M�UW#�@���"(	}���5���Ζ�~�/���dan���[�&��$�Y�%���=��f�T{��u}�� �Q�SX�S3NWRp����2Ț��3���G�[�D=i��z����75���T��F ��:��w���85㢂n��g�_h�ۏ��m�4��#��F�u�>J�&�x6d� �-���QY��Y����?��/?�`��|�-�"�iuP\�elMA@#��y�������&���/�ߓ��E�=��<��]���j&�ZB�GB���p^OO�~DO �/%%%ɓs�0;/���M e{SX�cF/b����ւ��B�Y*"**�Is�ޔй)����ၫ�s���6T�3~b�� n��_�G��N],Ėc�9��!іd�V@���>}�l�2u-��S�+���져�|�L!�����)�r�{zJe�x�;�7�<�Ig.�^Sb��␄8���F��q���h�ԭ������k�95� �S�11��Ȃ�@�k����LϿ��z�-]��MK���/�!$��������FAK�A-9eC���N��s�\��x�[j�s��A��{�6�� KB(N�SI̤�^p�'�?DS{{;V/�H*"�@�JC6u�?�6*I�9.��]Z��<kj�2j���͛'�a���F����,��o:f�p���\�
J���&M�uc}�<���R�-)i�8H��AW�A:�:�����Ɍt�*(ෞ����~|�J >:��6��ņ�ed���܉Ȋ�+yu��*C-�/C��?L�j͔��{	����r�^ ��k(7�4��$V=�	�U��ng��x�@qܤc�;���_�*�jkU��*jĐ������&L!�� )]��$+�E�?������p>�_]�p�����d���hˏ�]��㸮`��"u�����It��
���i��y8���f{�={���7$)���� 1Rx;B�6T[E�?Խ����STYY��8��i���kvv��^8��n��0X1��[�註�ɓ��H�ߒ6i.jř|6��5G�ʳ7/�OB��)�vv��ĩ���Y6�Kq������kɝ���p{944�:>>��q
�,Ζ4}�=cF��l���c��2Nx�������)������c%h���J�tj:Xt���^�s���� �3���>cFRYC��EM�hsNk~o=�M��RK�����"꨻:q�Zhd�_D�$vU�vu��
�-����dƜ�9��ܩ`c|g�P����:ܱ�����v݌2��@�(�;�R�[���}E;e���BB�ׯ�lE�!P���H2t���+�f�+��4*��胢�r�AH��������
s\��#,2kٲe-Ǖ����d�C��-	�v��t�רm���(	Md:T���čj����:w��T"��>n�JK-na�T��fM<�X��%,�V� ����iOi!�ˍ
�0����-B	d\�3��LF����1��G�\��eu`%����B�����.�P�M��8KV	]L�t�vnAa~����F��� �(��ʧn#䍠�,�~(R�=���fc��������"&�e��*��䯽T:�|l�+�*}98�h,z��Fc�*��E�;J~$N���[ϑ�-���f$u+,2�c�Us�m������P�Z~&y;�H������>��d	��ɘ��I�,C�QUPQ1DwlS�.S�����W[m��t�����I�f���Ѝ�j4fs�����86�v��딅E���F��`Km>|�ø�ĸ�A��u����d��Ý��;���b H���%]I�~`�)��,newi�Һ�e���~.Vl�NQG��� �R���n�����a'���DP���PE���� �&漁�???�-^T(>�#�uQ����;af�9�F����J��0&�:�!`~](�Ѹ;�Z,�e�>��m4�Z�`@:,3ĉ�j����P���� ���
��0Fe�??�I��j�o�����.��r��-,?����i���Q�n���|��.
rT���u�0�y����$h��ʔ�]��X����`��S�U��pm�S�P�� �hHS� �(�ni>���ゃa!���mSb���8�oKS���V��h�|��g�I-��dS�YJ-�������|F�����W����}q�f��uA`�S �A�������=�+9�2��`���F�F�����}H���H�ڈ���[Z>N���\��X!tQ3����ͱ��/씱
g\�-?�]RR�0�9�f�P���n� /��o�@9�~jRC-���0��F�E��F��<�e)Yp}��3NǺ�x�������f�jx��m��F���N��l֨����@{
JJn�p2�>�AB���#���b\�a���Z�b�Y���N�]�J��j�Lvs�]���W8��')��;-�s�]�~������ҌWb3��7t��y�A���r).��Z�mgt���$@�CЏ��{�pRL���!(555�������
�E��'�_��t���(�ۻwo����_H`��dd���h�q�f4���`��2gv��r`n?�Nof�s�љ�ϫ@G �W��N}�1ണ�cjr2�G\�ǣ��3���J����c�ݨ����JR�JY�7"ԸC?�ΏE)�9.�����\�����G�������e,5G���~*�M��CU� �
_gq^��E:)���w�Jbu�bG������ Nd�}�*��P.��>�4x�d"/��.�A1��F�V����W2~*#�E�E'G}H��<h�f�����d�k���erB��w�z�3e����e�{����}������p3�L���XRJ�WWYT�4w��|/�.����c�GL8t��h';� f//���˾rT���<qpwA�7r�����g��,��۱�����H�rRr��\=��0�1?�@L�����o�g5G����o�z��n͓��P ��W�but�Y9KT"K[<������S��#��������v�������>P,�� �78������s4�eTʍ�_m���,�_9G6t_΃���#��s �wU'z;2Rt��Hڛ��%$��֔3q�3���k��mB�}�l$B����K$���&��� �nnn�x��n�OhM���p�g��+W��%W�b�{r*G�#��S1{���[��w�U�┉���Q�эS�d���	0����?����P���H���G���P�&'�����Y46�?���,���.f��S1�@�����IM�y2T��b���@Y06�}R��ɓm1B��q9F���#�;�er�9�a����w˪݇CӘ
��C��1�l�N<;-�i��U��%���`����^^#sdM� �B Ta�s�����IU߂���<5o55I	�s���/��֠�F|�\��G��w�Śs(u���1%�I�'�F����	�(ऱ���`�J��P�Yvu�;|���	C+u͕5%߾Y��~i�@�!��# �L'�i��=������G��3Ô�jao�U>���S{���s.u��Mʺ�~�3Ф#��
���ohhPp�)-8�8���b���MT���ԥ����@������(��kMv��;枃��� ����a�Z��5�2�Y�zU��޼�Vi��P�37�[#e����9���L[�#�d�ɐ��S�ټ;���Y�c�����n2�"�� |�N����":RJ��p�Z�����_<{�i6k��ʷMv�R��8�8i b瞢Yk�x��
�b������Lf�=����,�_�?� d��k30�t����DmIKo��ĕ@#)����minc�㋠��N��P[H"�')Jk���L�	�bpP嫑p��1�oі�ѭ��wO��ߌ	C����������u�WJ؎���+u偑��Ē,vN�6\o��N5">����T������w6g�D~��Uw�טn�-���l��$Q�BX����.��(��luhv͊�oy
���Lg[a"�@�
�F�eg]�=�������1SH�Dtrtt�̃!�٪�*����-��E�����g6�N����\Y�#�g�:�!�RF����!�lLLLSY����m�;��"/o�u����������6������!PM�����H��<wvvVXF�kn�N�e��#����iH#���
Q���Q�ub2�:�
���3gC��a琒���ɭ��c���n���Q��bo`��m6��7�5Y�2,�N�
*H<��ġ[[��	O5l%6F+��}��U�N\�5�9K
����,��A�Ȯo
5D��x��0����k[�3�5@�q��\A�T���c�;P\}oP8 şξ�2#4%���(b�&�d�^'�P��i�L��
m?ť����-a%�iFH�?�� ��[�1�K��y����<�*,4t�G��N3��X]]]�@�Z�qR\������O�*_��n�ƞ���]��3��
]���ݨ�1�RI]��d��?}�*-)y�␻!0��3�N�U2�c#����Z�s	&9!׮]���	�C����s��ul�*���ɬ*�-��8����u˚��ZXvǾ:(�s����<1q��O��.gZZ�e���7�(~T~�qwԇ�sO�n���p<�>���(���q:�^c���ju�|n�FP�J��/���f<o*J�˶J����8:9�*|��BI�k�-1�p��0�Z�U��"Q#U�wGݠ�Z�ӈ~�m|x��*mL~�LG\��d���01.H��O�F�s[���~��VosW����i��|(���)�^�`��]�I�|x�]���szhx8����vŤ,�|w	mN�P����#p1�ݎ⪟v;�9νh�>|(���S�f�.q���zFF�>��F��H�&�r��O0S�� ���?}Z����۶m�ɰ����Ay�����f+�b��I��t�d)5:�� j���HQ��7� P0r�j��ǳ1Ϗb�׽*?�l��+d=ř2QlNA�:C����IV���qɞ?����)�?G_*�2]��<)�>�T��"�����U8[Ҽr��&�~S�a�w���u*pa�sNYD)���@�N�8�`啼�]��;g�-���^o�o��J rA|��K=P(0�U[���K�ۊ8�(S���'~�8%7\n�}��Y���R�0cU�ћ ǀq���ޭ�o�b=P[Gg�)��z���iiU	(W-���
i*�)��*����肂���U4�riiitC�xdVF�9ɽ��2+>7(�ڟu�c���]:uo6��x�ړ}c��o
6ų�[l�ɼ�|�w#�O7�/N\���xl8�|��ݛ��8������2�w���B�+V�)�M_�h���d/t_�(~������/_�|���;��x�L�;IjLl#���,}���;���MsR�tx:T��cN㥆�4��!>��}9d�c��)4?CΫtp_�n�JK�v��ƪ۶�k�%�U�.l��cF�3���vySs�/������nm�B�ۍ�eѝ�sr�V�}D������P�S�c�;G�ٜ���.o��~}�a$5fJnl:��ľ�z���W��]��۷:����Aj��j�W�����"y�ګg�B��i�9(�G���;����
a|{��!����o�������w�÷���u&����Zf9l��K��:7Z����[k��>�\ڄ1݅��ͷ��ހ�_�y'�}r�s����d��&2��@e�M��99���~5��ֽ}>6��oP��.5�	#��
���>�,�qv��<� ��3�U4��_fd��{[K�q]%�l`|��q��xX2��PoKR��,d�s&FF�I�S��m�@����aٹ��*����v��7�p�4'�=�|*b��cVR���Z���c�߾=	�9�A�@Z�,
�55߽{���uF	��ú_�\{������\{h����Ȉ���䋠ht�)�u�_3z=sTSr�����8���KS�g�svK����t��܀������!f��Qf ���y{_���ŋ��7\R���:�h8�|�ңŤ��<6�)<V�A�j�:e�r�	��~��e�aO�}$q�n��K��e]���#�ء�)�d�>D��D�G����IS �i��v'����a�z�PZ��QIA?�T��Ҡ%��w77�F�� 7�<������J�𲉿�a����`��d.��I&��K-�CG��d�M���N�={6fS����.�?���-If,��b������3��[-Q�$�Ӯ"l�KY�Cv�YY�J �_��j�"/��"��2�c��q	��wa���V��\��2	2L��6^���,&Iu��/������R�,N�O6b�ݦ�(���B�w���@��\l�J��f���Gƞ�.�����F1r���w�ܴx~�ڭޜc��taQQ'
��>��]㿀���@�-��O�Υ�����mD��V��o���S��c�B�̊�CSU�%%�$ �3rK��\�e����ߤ�Q3.�3jk>�60���%����}�;�ī�.DBo;�R�� �]RUq�rµ�ĩ��9��j����A�O]��'��J����0^�����2�2�+MvK@@8)�_�o�+!C�ގ�ᶸ�ޖR�HGo�-}�Tx��27���b/SRT'�rr�a�sw�Y⿛�8�4~Ǣ�oUI���ሓ����9��§�5�2�X �q�@���|FqW���(�yvuu�"{u��؛U��So��!��FJu� ��c�`��ħ�x���%/��0�܍��<x�`5�KC��杕[�Ғ�	{���������u��x�!_~�Ҏ+�4��U�sqI�k�P�$�3�CK ����}A�:��ó\?����գ*�+ �Nɬ�5�4coj{����|����8��CME����y0��A�JI���s�'�d��HI^^��#2wx�&;#A��zkC����2:R��]�I�|�ͨ��
��9}h�=aTϽ�7ⴃ��S�晑T��·1GpHt���1�m�>��[���G9��n�[e�<�� �q[�$�b%�d�޽���G���6�<H⤤8-:Y�m�Ɵ���&����q=�3J�SY�\���^���,�W
������I���
�	��\r�D���j�Ԍ��m�y��%$$�as��3:im�*�� <B2555姰=דz�������}�d�A|$0�c����~���e�ov�b��A�P8��4У~�(��2V-}���U��4�����'��*D�wp	�	 #Z�`�A��J����:�Pj����8ݠ���R�ۥ-d?�n�����nn#�E���a������p�ӄ?��}��m9UI�JJJeX(��X��ء&�ii[�Y��/8WX�ϝn9�W�\\}3��:{(zjrm�/S��ñedd��1�H���H�����TfM'Y�&f2}uu%C�[Fa$ �����N[��K�9�� '�(`6֟#�`�el���k�C$��5����dK��7��<�4@*�nR�v�^�����,�:����sa��j�-	�.��7ߎ���Ɣ�C�ݴ�K�X�!����	{��/�(�2�F�M�';7�S�&���26�7X�'��Jnnn��Ҵ̨�SD�	��訨���(�"i�Y���QE�k�=��ɺ��bbأ����(qY[[�'���d�j�vO&3�4��������b�!�8�b82DI�I�����S�֑���m�NF8�sv:+?m�u�L7z{�����0���D�$��pz�%Tj8!�)��ۓjg�υ���k�Ki))nz�D?����zl]<���M�	�XNS�R���d(�B�_��^wش��L�M�;$�����'r�{�p�ǀ���?cR�'�*��<�K%ۺ��[�(y�@���t��0��<גl����5'�����w�H�_cc#]?$-/{/[Q[[;L�)PwW 7�viW��Y��[i⵭��gT��:�A��/o�O�H�UA����	I?E������P���GZT´Q��V���(��W�Ț]F�'KSI�[�ƒ�����aJ��
�G��ނ~���9�����/�}����<���,�s�����̍���L��p��4�z����v��_�	Q��۫����_���� ;�{�s]J"��[+pwj�@\Q����x��ͷ��x��D���+o�ǿ���[.x��(�yak�1{O����(5־{`��1^���*�w`�ث��B*n��S+�w����$�OَʀΊ�I�-��������OlVB͉'w���ɚ���G/�2�����7G�#b�� ��g7�|N	(o�f#|B�x�dS5�lq�"��l���^"�ߒ}���G׭[���߭�b=y�u?� �4W(�O�nĳ�_ޯE�ree�E3�#k�M��d[��x�/�0��<`�4�^pkkkJZZ�	�BEQ��PR:�M�v�?z�A_W26𗯸�k�XK��O�>���=Y�q���(7�X���9�.�Q�NB�9E轛{"��Ӱ���\Ł>Cu;�㨑d�/��8�n)�0�U�W&Q(�F<�d�nR�$�
nfs��4����M���]]��� 4<��7��0PR+A�D�Q`�P.���Z2n�a�6^^^9����a�#����^�"����ߛs��3l����ب5ۼ�_�!���y�ga� � �~�b��4^��]%f��Ñv�n^�PD��.Ĝ���/J�����rq��c��Q�jR>I��A�+�mn	{z<�b��~d�b���X��]������ؽXzV������z�� d/�]��&�!����5�p�s�zn��U����'6�B�@�|�)h����p���+Zt���aX�nb�lsWD���-"��R���v�qb�V� ��v�?%;(���e�l��rA��Zy^ ���Cw��bܨ2	�f��f�"�~��Ͷ��)��+�I���{�����aL�Pn�O�6�s<(�Kł��kp�f�����v�oOyd[IP;��l�=۵1�M�¶u3��(	3.o=)t�#>��< �S�T�y��k���d�u&S�%�qHd/�n}������0�\�������瑧��*�e�B�.!�b��ح��?{^�5�T�����ͻb�y� }��É�Y؆��7���ěA�O�1��lq#B=��u�u����؅�3�=�Z���PUK4�]{�ڶm�7E�Q�r�XX��]x7`	e��G�5���5~+�e�
)l��^g�g"zI�Ph*�� ȟo�Z&(��p,�y���-h�孕3�psN����W4h������Ӎ.�Q�|�q#�3�>�X����"4=���<#(`D�������I��\��f<Oj�	E}�M��2	�5QUchV�-�VB�2G��ٚ5��~붉���~iI*�������`m�al�bD�-B���)w@f5Z�<�s)re�Xd�����V^�t/Gbב2�CO��7�F��6w���z^��
X8�*CU��CQ�z�A�]��>5!����铃W��F��"�~pJF�r$���ʾ�r�-Z��[v#�	��5=����
�=C��ODZᰤ��T�ķO�V��l��"�d+A_NBOV|��9�1c��{��En�=l�`j�g�A�/�rs���+�x	�^�GL��=x4Y ���/~RD[�эj�;�Q�ȝx&a�s?� ��D^�{%������� j���{L�<<bjU:��N��"{��M��������In`�cUUUx����^[[���H��ߔ�F�}$x%�{d؅˴���pD_��(�y�˯_�ЍS+� -���qy/
C�H�[��63�mnn��k�F��y�D�P_n;jR-�'��
� �ݸ;�yH�c�E#S�L�/<4��o1'��<y�2Q��C@
���M��0A��M6����F*"z|(��0X�p�r;b��8�yب�]�ty���M��
ٌz�G]H:��<>�H�&l�sIlZ�,��J��sm�q�,��7�ܪ�Y~�cj���`�{?�$���iy�,7�+~A!�0*%�e.6O��z��tLsGu��ː���Ti|���>�9}����rS�O.�l6)/����[�+ ��}�8m�]��xIA�K}��]�F�D�������(��h�'ZͫFPs|�"H>�Z�X���q�8Y>uC������C���(h�K�i�㘺��+���l?r;�>�P��$���+����;���]��������E%���]1|�}�T%�)ytd�l���/��C&t�&\.%�WM%�9׽@�ElS`���䖍>l�`��8l.$���ͩg���bc���Ԓ=Ӫ���G��`��-1(��T;:kh�M�� mT�i$�ȶ"�uu���&괪��l�x(co�d`��bȍ�Z�����|��`�?''��S�.c�4�\��1V��o�C��|�;s	e��IQY�x�����{� ��;���*��m�հ�sswI����f�C�[�9���+$�ʮ�V�ݺAA�0�q˘����,ǚt뢓߷"z}��ωcM{2z<*�ܭy����ȃ.��crjMTi���	O�v.�Gl�z��.���Z �w�WB�0�Kt���mgV�A�VF5ц���2	t<l�oA��Fnk:Wz��4[�o��F=D�͋�j.��a�=�ͥ��^W �s=��)z����!Yf�x>K:X>���D܎���P-}V��M�nz�J��eۅ����-AGQ'��Q��;g��o�v�Z ����ڸ�ǈk`�m�eQ��9�8e
w�)���^�F|�
��7s j__.�,�p�w'�����/i1D�I���̴���A(k�:��$�މ�D�Jx�sNl:���l���q�<tw��fQQ��Ρ�HT���=�sY���U�=f1���-���i�^��f���K�zNd�ǎ����62J����w���λ?$��Z[[�U��$#?����bS+H��?��3y� �d��d�qww���5�ޡ�-��2��@���#�5*Y�-~+�&ê(����phc�Ygo�>���B�Y�����5�(6١�
!@���x�Q���6��ˇ��ՉoI�u�w�ō��d�=�*v{$��B��h`� �1G���~Xo�_�˹�J��)���$�з^m6���`�]�ws�U��`�Q��\׍C���+sh��t��W���4Aa	����}�3@Y�~���zJ��4m���z<���)S��^ے}j>�Sa��YA>�s�ώ���R*��`���_�~����#��ΐcT0�"_籐����Hn�*���늖hH_Q��T��>z"�s��-S!!��QZ��4����������]B��Ԥ������3���=�-�������	b���á�
D�	�������@�Y� �5طg�Ac��f�U��x8�n�y��j%hFY�+ƞ�y8>0}kLOa3�P-��LP#S�3�8�;�*UR������)�rP���;� F�w�3���y2"�3��WG\�y3�����@y�P;ޕ��Xt�7&m�������N��"�a�}�C!��s��Bz�V��ړkQ?����1Q���OsA!�d3
_��*�&�ay+�V�@j�q�w9��E�.\�
X��/i�g�\ga~��c!�_�_�[�Ե%��������|�/E��)�[\u�1O�!k|�=�gI�����w�G�V6��555E�YQ�ZW:���qcwH���[_Ծt�v�"D���|�u6���?���N��!�"
����EW���A�}�{э	{���<R��th�� C�g`q0�6�I���&��h$~X(��7xi��}j����uttl���{f�ֲ�j�������$ԧ&��B	�I	�/�֓�>T;�a����ﴥ��jk�98?9Mi���	���{����5�}ſ<���8�m>���gyܲ(X��B�i	{Y/�!f��ϲ5G��wT�j�cE��=�n7Bf���[�94�����%,zt� �u�c����ϟ��v�X�����l�t0���誮��O�IAq��s����DeQҘ/}���h�(1�h��g���\�աR
@�:�DMd�o�@|���ؚ���3s
��\#��j`u�͏�6O~~���dSK�/w�\Ɉ^K����Yk���_�G���n�r��Pֽ��}f:#�<-�kW�(g�呁v�vH� �D���J�H��UE��u�5�M�����$ ��d4���$�c���$T�µ��k��7�t{�',��X>��Bs�A<�nY�������IJO'52C?+�C�i������v�/���t4���n%C��q�	֟K�c�褭<v��$�� ���(�݃���/.��)���zg^18ZQ��=�S#'����Z�4�s���k��$I��{Lq��8�C��z*�h_ߖ<��5�{<��]�*�؅/�sL3��,z��WJ��gc%OZ]א��&��"���\"��w�d1�PF��4�ou��	�������P �ʇx3��i�V�w-B�����.!�U#b��(������6QN�~�¹���Ѡ�V�� [�Ѿ�zw��k!�X�$��b��N�PaL��쉢��;�{Pz�r ��>��;lb�e�v	IC��~sL������OtjN���<�T�7:����浕�NCA~c�~Mь�?{�o�l�ӘAEC
�;��J�<��y�0����V��X;��_��}�2$8�`{��8q2����w���L��7��
Qhc%�]GB�is$��W>\��� ���R����ѫH��-:"<�`��%���+�m��r���C�M6��^�0ٚW��ϔI�F��Y�g%쏨�L���d��وi��5&��v_h����O�]��d|Muu:f�GҪ�א������Ʒo�y�N�"9���|�� �lR��ss`�����K=-Q���Y�:g�_woٽ�Tp�����+
�!����3b	m��:)��~fc`�`��'K���Bm{woQ��W\i�Ȋ���[��ͽ&ʥ:�����6��W�����4��;��e�ꛑ�}>%
A"/��uaL]�\Nm�*߼5����7o,���J�G�S"Y�����Ʌ1��2���z�C�E��\�iڸ�AUB�R�WP��=vS(�O�ݢ�5��� `����R��xr�����+�-g��<�&����c�h�[��Ѿ����g�
��X��p�:�+��v`D����
�S�ACeeecG�\<f�lQ��'�\���	R�{��+��oT��ن+�6�S�_W��w�/	?xv���􈶪�Y*<6�.O}�0��cA�f�R�_�M�J� ��9}�xw�������F���)��M��-@��4ukM�yd�H�w}o��p��[�����r�����w��6���,}=U��j�s;m���00������o1��
��M��aN�(�ns������Evo��^�*`����~++�����G"#�	c^$g�4|�P�^�W����V���!��n{_�c�]|8h8K&A"�T�	�1T&n����Qϊ��ʗI0%���k�RL��G��R������� �Z����nm�,w�a�3Ӌ��*�/���r�9���&�gL����&�tx�ܸ<��e�����<��2i(A�q�Q�D�衙�YײXm�sk>Vǩ�&W����q��Jl]E�o:���;~R�H�IE�Z�B`�6��J,�+���P}:όG�BcZ:�<r-̇(sY{P<DMvN�"E�R5�+��XE�����E����=ܻB?�t�U��0�p�`�h�h+w��.S�OG��ey9�뾚���<߁���~�
�!s,����(D�l"�=��Zg��=���
���G�3p��?@Ku����Rj���=_����^����L�8��k��^��i��/�Hw��(98я�G�t��
�|@�w��X@����s\�s�2/8R!QΨz��r��*	$ް�lM��ޚX����mn�c�Ѥ�O[��n��|ི���L=)p�����Z�-ᝣ7�~�:p��]��:��B����&�W}�;;]��R�Ie�xc�&�"��f*���lח�K"��[�U�C�t��{\��g�MGF�t��I��Z&�¥�|
[K�Ъ��x���K	9><���괟���P�d��y�����7*`
o��!ڷ�z̠P\�'�*�n�(�q���U*d��2���V�$��`c��3;�Wƞ���>f��z�p��n�b�E�j�O~��!��d��y�GW����}�St?-�j���u��_��̑���1�2I>����^ϓ>��*�J���]��d"���[��W�V?Z�Q>v~�Ґ��澚z��aa���>�
�:;��������Z[�k3����T;C'g��GcY�\E���1tsd�{	Ꝕe<�a��4+��e�|��-l�~�c�E����9(/�ۦYSZ��D��TE����X,�&�k,]�%>h��G��e���S�*1U5z���HcX�6P�u�v���T��]aU�q�4�,�-l���|�0��^־�7��~zW��{��ٍ.m��<�>�X>ͣ�j'k�*D���aG+�-u���&>��8�Gs���=�bt{k�4-��խ}����������B�x�c\
��9�iU�4��H�n���@]�=�N�h�5ED�����T��.�B��Nf[B�_^�kFPy��V�G������G�m������X'�Fcxa�}́�"�9�̺�Ci���(������s�Ѿ_���e,K�;�t�	�|% ��c�ij�*�cYn�n��*��\6��Y�k�UOKɤe58Ǘ����pVVV��W-"��#:21�{�v�dk�j���HgK"f�_��	��̶�����Vd��Zt���C�PA��1�|n���cc�49�\�kc!n� �i��K��b_�zf:��%D����iT���,�χ,���LB)��|J��<�pH�r\�	����8,�����x��H��Y�#!����A���g�L0ݩ;�.w�ws%b��6�����Bz<@O�H$	�c��yHp�]���hk��ЧbW�qow!��:�'r#�S�����p7�Myw4�1]ey1����j�鉪�K�i�FM#����i���=��8,i5�%�����kac�ϊ�h� ����ސ*1��_� �s�b���4M�Y��s���9�����ZK-o���P y�C��B	e{$�r����Q�'�E��l%n���8"��X�bUaв��[)�1��#亃��J8��d�P�J�S62w+������6V#��v\3r���ۅA�+R�.Yn/U���飏Wz�¸�o�%� ƹŬ�e^�]&���=��EV�
��i�j�c�$ �t�n�>�+X��ȿ� ׇ��,ӌ�	.Ó�G�0��J��!6t@�o@���A_��P�QOXE$kk�%ƒ��I�>���J.�MoszW�I!����:
d��m�v�r��$�a#6U�^L��y~q��xGEE���;��H�K{�1?{71�Cl���t�3p���T�.0_o��8&/�K?9������Ǉ��Ch�m�R�T���	���f_���lꝖ"���Ȏ�J��l�=�P$��-�����]�^��)��K5Q��8��w|x܄�R(�߸�@NJ�*���.I5��C�����o 5����k�Bs��H�=:2���	�:?���$���l���*F�D�&ʴ`���ÎR�c��<D� �-��[n��o��0��"p�_��1aaa֩�[�G�e��"S���u�
����+v?���}cIv]�V��["��U����ׁ%�d	
��A0m��Ph˾����i	�=m�����'�s�p�~@/b��)}U�� ����K��&K���*'i�q�.ʠ	 %n����������gʺ1B���{��U��L���^ z�ZeWd	�b{��`8�³W�l�Nt���?()C.��c����Jqs��+�}Q(��bbs8`jB��|g��P(��3n�r�A]T�)���$�I��".��"�|ZJ�s��]���E:�O�і�tT�Q�t�gx��.�Î�6��1�i���m�;����q�X�$��sQ�p�`���OGF��s�([�	�:7�ֈ�~] ��ĥ���v�����⟜�[C�Z4���X�/�T�J�+|0�޸[���Įԅ1!���Uօ�A)ѭB��EjXt֩�����-�W�g?�У�Ix��=EW�^u+����c?�%X��xB���IbQ����{�*�fi�fK#���GGG����X��WB�~WA��W�:��&ƜU��
@4����?Do�%���i������ɡ����.ז=�s�NT�
$?�L���n������w>��pOF��J1Ns��nb���9q�PfK�r*�aǋ*ҩV�#ցPt!UX\�SRbt��3���3�M$�L�n��
X10�����Ę���#� ڣ7��q�O��z#��߼R�[���<�T����5~�뚙6ڊ^�	����.h��z�VT�4�6<�e����g��nӿ���/\�rh�C���W��^r�����6��@e� ���B�D6c�z�0��(
Y�
���� pݬf/����Ry�a9�tr5c��>CJ���`o�6�ȐU?v�IL�Y��D�-A�&=WD� M��Q�pU)r�{�{

!��#�;���[7dN���mX��S�A�H��r���}Aľh!����
�;K�4���~2��	9��N7Q�vD>t����g�ea>�!�Έ��E'~"�x�>h��,u�h(1*ڂ3#�x^�r6�u�0�'�U��{�4�)"�Qߝ�tk��H��W_����� ֓�5�U��g��K�+�_4c���_�Ah�(1�V'��]UG��}����&!�gS��N<���@/��І���R���b��S��aJ��"�h�M�[`�6�s�*�{V$Je����tH�Җ	dC2dT��cnj�2���8�H��os���x�$�9GN��Kl��𢡊B���C��R �x��0׃�4F��u�)���mH�~��e��m��|�y��	�*��>YFF+�6>H��-��N�/����~+$ǵ��x��f��Py�ڏi�5ȄBTr�t�.�p@1� l�NY����\�9�'�h��m�22^�u�y�U�^��*D<.�6�\�Q���c�i�<��&x�Ω��gMT��\�p�V# ��;L_AQ��؎�4�C�5j�K}���U����=;�A��H��+���T����v���>�gBm+J����^�d�ᎇ�������.·���`�}��#��m�M(��92�"\,;K逎�!��̙�'�k�I�׻5Fn��bTݲ��D��"�iz���z�L�-�9�rfF����~�
�S�<b����=��Z��<�4�T����[�-���DT�3B(����K��.m����|�\
j����0�\`��t�������C�Aa��>�+�6/��,4^�����*��� ���}��}d;&�����xJ�ء.-�sx�.B��N(�~#U�>���}�a}���x�7g"Bh���+S&��P�Χa�{�\�w#۬A����Xc[����X445'O���>:��j�4h�A�D]J�E�	=%ƅ��t�{D��]m`W<_��K|��-�<�I�u*��.1�C��)x�Ia���Ȝ��Bn^�6`�je�x�N��r;���\����"�	�1��_�⓵�kZ4?!".S��
L��h3D�⓬TcbD)��N�YY�"Q<�D��AwM��A2j���J7eKbX$"ǋ��Ί�>�D��V�v���(=���d�P���o�նP^��ߘ��zd\�⏅���n���^�6����緺if�Y��,�/5M$̭|S�.�V�<�H^ؐKd��c�hր��c��((s� \��S�EWƌGi��7H����FP���]�Z��Hc,J!c���WD�y�nm�X���o*E��6LH� ����]u�qˑN�5=�i��'����Z��w	φ|��
oK8�v�$�[��7�_��C��2�;Q[u�
i�	8<����b���ⲝ���Q��v�n9�6�K(��\>���(���Ǭ������;h�ӡT��00�[<�t.�C�P�s�l�ǀ�(��.;��.�.ׂ�f��P��F�_K,a�W���Z����gx;����3�O-!Rl�ݑ��@X�k��L7���Sj��:^"W<�.��A_oŬM���u�S_���I�E{�vI�IyI�����3�I�C��.�-H��R'��/��誧>猎�J�f�ڌ��X�|�)ڛjb&�"�zJǼ�Tm��8"�$6{��E�g$�a___7h1(� Em~�6Qlh�-\v��ǌ��� �ֹ�!n@0��D����B��Rï�0�Z� 34�+J4q�.��s���GjJ���7��6�`}�Ay�>���	;�����^�ʶ��%��bE��&��p�|����J����r�|�܁�*^)We6�!� W��i�S���������/ ��9���I��:���:E� cu=�}�2�;E7��2��/8��PTB_���r)@[����y/����H�vA�6�u��8GnБ�$�5,=m��� ��P�M|��܋�a>��ȗ�d��`!�
���i+�C����z���!���>������R���Ĉ�e	��e,���Q��@\\\Q
�N, .LI���r5ǒ�?h�N����/?�6�5�������glb��p� pp`��;� ��~Ӓ)��/k՜�I���\4J1+��t�>���->C�6�x��qq�3qy�ձ,�GP�Ğ�/?}F䳔O����赎Od��>P>��p�d�E�-i"��t��W��D��7q3sWL��4�
J����S���H0�Y�����RL�FzĻz��P�9�-Xh��sҷ2�L�a}��r$��(����o@�t$:}vVe��v3��̚$����6wn�Z#�Us�����S��bz9�b��rԉ]H�`^C�������n�I\� ez��
����Es���E��3�Ǐ����I��nb�1(��'�W�:4�Q���2��5��5(W5����}���K�	�gn�"ӡ���gj�f
�rW;���ئXˎ+)����@]{�>I�=a=oh��sà��~���D���k�Q��et�&��'M�����ܷHj��߼Ÿ�7�z
�qLIŜV�8��d��f�F����!/�'�v�x�0�9V:�n�0�(y���(R��N_z��i�:7qziV�Eņ;E�D���F�SP���)g���(y�O��ys���;Ґ�= 3��V�a�����26is�J�11ty�٪�NvNl�S��w�	eV����J4x[[������Q�kj[D���}B��T�^v���Z����f�_i{%:�dj�(���,T��D*c�n�{�Vs ��߀s�q& �ɻS:�*��B��iuy_�!3r���Շ��_�^rqZV$+Ж\����7un��M ��@�����E��G��VhE[��-�q\VQ�=[EE���I���������4�d�i�|
ǯ E�sp"M*LzXn6��l߄l�_4��Li��.0�'��_,;�<��7z�ƚ�{�"�f}rFg��F'�/~��" }w��>-%�Y�慽u�9�A����6<�� k~o$/c�:t�@Y��zеԏ5ۉ˪���R]�ۍ�����[�l<I\t{٨V��{3.n��"8���"�d�Q���������$�4��)����%�)��i��z���Y���ϯb�4���+��I���k�JWĺ/p
�X��m��>���3s�XdY��s�"���xן������/��ײ�b律ⴵ&� ��ZB[��_7[��ˉ�'���Q??��������d/(�u�,{{���R�(BHӽaB^GN.�T�������-X�P����Ai���0��6�D�ӭG�dH~�Lfʇ%J��䛬D����`��`�KVQ�w��;��|y�������L�u��1�9��P��P������䀹i[���-s��S����I��������y���C��e.K�tkϓ#"��.�՜O�x���I����]��KPbӜ���#GrCo��.��@�H�~\cZ�� *)Ɩ,��-����^���:sI؟q�UQ��d
�V/�����c�M�V�tc������jv�}��r_�c��Vp��ag�-C�&%?낌�2ΞQחQ4|BD?F�s��ζY.���K?�x��~�$	�MZ�I˧?�I�Fm��y�����Ͷ-�z����\l/�ԁj�J���7�jS�7��_C�F��4�d��֒!��ۜ]?�������|J�5w��A��Ľ���nH 4��/3������ ���	h?/�X?��q�y[�g1�s���+�b���\��R]� �p�_3S4�����|�`��6Y�/�Vp�K��~d+�]O����'�|�VW�d����=×�DU����>G
Y��d�tYsb�I	�OO�V�I4B1�QJ�"߂����}�)����� ��b!����1�/v��"4�3T����dn�7`��"T��kj��ͧ�6dY�V�N�鿇(h�Z���a��P�#���N{��&�X��lL̝�izw��^���g�т5I]���r)P���j�EJ�{8q���O��{���i�Ґ��Ldg�L�!��z9���3I�S�͡�!�Lm���+�V��C��/�zsǩ��H�n���xr��W�44�Ox!���c���P�4�7w�N0�	բ����l#�?��+�[�]������r�:HVXۮ'q��j��#�:���F�����Q�ݽ��g.���8�~)i�Mԅ���{.Od�	�F��ͮ/�� $�
��Z����Cd����I��v�՘�d�P.Rq�n`�����9y���-b!���L�Q2�𬍫7��z�&XL�lҢ���͛-j-s��TfNaaaZ��?]���\�;��VZ����=\��b@d��[���[��O{6p&�3|DJ�$��'C���o��c�8��E\�*-j�}ٶ^�7�)Z�k:�]��G�"{�bּR�6]�w�%�e�F@�~��ږ#�k={e^{��M佃�]�O��b��ݍ���G���xKP����]e�n?�D�v�J-�G*��H޿���C�'��	��F�&kE�wT���5�Q��ӱ�]�Hjz6�<6�ҁHT[/0;�5'����')�i3�ޛDQ��0���i ���"�p��\R�ս1��=a,#�eVw���+�ߑE�U7)�6�Ns.�1M���y��&g�ScHݟxm^�v"�囧c����1�W_�;q���I7�秤 �e�0�. ��!��̀,Ϩo/()�<��o�@$u5��e�=�L��[������3��"������5��hTD���T���[�#���b��R.�6�}����܇C�d*���y2�S�f�b}��F^��g&�_Ify�\���Ə��b�a/(��͏�m�3X�qN��h��w�9?�z+r��$�T�l�&y��ȘP�`ˎ�#�7�Uo�����^��Z= �3�%�ۥ��ѣ�T�H�;��~�M0���?gL���#I5mK�
�h}�c��+�ε�w/������kg��'��h@����h�VE��jW�B���X*9���6̹�^�E^]�GMH5�k���r�<Sg�BRS����\>V5� =������͊���͙
�%�S��������y��EÚ�����4<îs^�sB�;�O]b�i��#����tΌ$կn�����Z��8�39C��\1QrV�F�&���(�D5�	F�̇�{<�I@luK{��RpD���d�C(m��1@��jD5�zq!��q�
wD�~,]U�+���w~Ո�R{�9jο3�3F^�G��_��S	�׌<�T��_*�9W1ƍK�t�l#.���3�%S���]���äΥϳtJ��+�ڟ�fA�9��.��ƶ=�X��a[��b�0��.��1icZv�=4'U��,�&MΪ�\5�����T$iX��齦�II^~�:��	��?�4����������n�܎�JY狐���E������ ��'�_m�)ɓ_�@�&��!��A�w����Zh�m�TzB)\J'EL�*-k"'��ɽ�������kH���(���j���<�'mZ0\oh���?��lI4�����s��&p�O�K�鄅|aW_~�:$�B��=Yfz��c�W{�z&(�݃\妡���c��v�֘��HA�M�E���݊JI��ʧp��f �C��j�z��GoN0��$y���2e_���w�r_(�:�`M���^~��q��u|u�����.���2�;d�v8���D: ��\| pV�x�=qm���'[[�LC��E�Y�ԓ�����9WI�������|�������1��Qf�}�s�1�M��W�B~��n����y��>O�W��{c�h��f"���"=�$U�J��76=`�ѱ�^^<���7���K�jo��p��N���@j_%��R/a����ݤ:�w��=y�ş��;�-��h�F�0��� ^^=i�W� <��_OZlE����Ɠz�o�ym����ɚ�X�o�o�U�u:�E��*�j����2���[v������h&Y�br;}�K��a�?�.�F��F�<)��ꆚOUj�
�T��F`�G��b�X�'RIqX���䥟w���z������|�ΗG��� Vhc8-vo)Y��R�P�C� �Ԏ�����������Tְ�Z�ɢ��e=!,S|��g��|5%��t��c�fr��(������9�?�*���dpKs�4��_R��F>��z|2�2Պ��ɾV���G�����!��m�:����0�C�򷏯���[��,-�W{��垭IQ��ꬨRM�D�wW��6�i����mq_�o[����\30`rt���.��"G��$��w6xl��&�������?a.�,Rk0���Z���)�r|�ț�H�"���5��C��̀��/?���l�GY�al�u?t�=4s��W���7����?B\��'%�D䔶�,$�Ψ��ۘ%��0�"�f�C�P<��~VG��F7������*��oE@��>M��q��R��mR���E\~�Q\ET���q�����`C���RSW���>S ͹#����<59z��#^�e���ڒ���2�SXJK"�6�9L��|=����hH��3�k��%���\^m�>Q��RF�&ҕդ���~?	!���k�?�H�(���/��x¿�mˋ;������ |o�U**���?>���A����nw�s\a���������f ��u�Tqc�����	0�U��Py��6F���Z���ړ�"��R�%�Q����׃���))� >��:��_����A2����n��u��E��|6�����f�.y�����E�ʿ�-�$=V\cmRJA:�U>x:�bɘ�\��UZ�T
ō��;� ޤ%ݸ�<���i*BR�bJ��-�'q���l]d*��;�5C[�D����$�C�ҁ+�o���&�0�1�M򿙙�b�!��8ȝ�_Sd5���^X���)���8���^K�k6����Yb�;7tU3o���Q��1�G����b�i�@��.Ss�`��*���f�B(����>�mX�8M��-r�����,�c6�}���*��MXwJ����9x��7�� � ��7j"�Ú���st��P*n9�B&6�)s8� ��ǧ��
�\]T�%�16f����S�7=����lT�L��h���m�y��ƩfΔ#��U�%�lip�)�S'���o��9��y�����)�z���0-ȥ�W)��[�ѷ2���9ØB!{��t*�HϺ$M��zu�Cv6��=֨����{��J�`c��f�,�'�u|o��6dFv;�y>�5 8�O�-���6=���؋������=�6Rn[#�R��ߥ��t���Ly���7v����=3�9�g��,]�@u4�d�t
��4�g?��K��
Ƚ����?|�P{�
DnD�� U*���0������!ޑX�֪�-�"�v�o�Sy{��B�p�fE��_��K*)����� hej�l���}t���:��j�]����C7��w ���@ͥ��Y fRf��3Mv�K�;[�M	c��6&O��4zaa-�%-��Ĕ^�B�?��N��<cH3�,���'ͼ �������u�b��pE\�����ƺ�����,���|�v�IGn"-xV+h�&�s�.�&Ś,t�B�������L��v@m���o���'��U�oN����~�*�����$}��@�:��7"#�v�����q4q��0.L!�ܖ���tNZ���YI|�̣�PԒ6�����w�}��ݚy�yC1�w/� mP�ܓ�;)��ܙ���t�ӫ���� <+�@�bm<��^sZ8{l('�,��sڧ�p����1a���Q)�踁�-*��K-��,��R��2��b�,h¬��`rAH	��[�ҙ���3�-8���	@߫
!�Q�uv�T����j����B�-�$l5�]GN�$����A���&=s���VD���)wܥ�8���q�;��X
��E����ωEĥ���@Mo!��m9I��1Y��$t�b�o�����E�M�al;P��C";���� U�C�:��|��pa�HB���0��FM=�l ����jF�u�uZ�,��vi���p�9��0�����%z�����4�3��`O��P��g��zL����Qt&�ET�Ĭ2TN*d�I��Y?��	�b!��ͭCW(�K�0��Z-�����~� ֲdyV�:����V(�|�%�~��V8��If�y����������S,�����`�����?M��~0��d$���a� ��4-�9y&���=4a�}N �(d������Nv�^����b�C���񎬟����������	�\���vkŜ������H�Ǆ�=�����~�9�Sh;�V��J����&j?_a��8�Ø�% E��(��`YP��B}L^�NEg&�nc�V��Q\m�R�ŷT���	���E�?����L�(�>L{���R��΄������+m�6���d��ɦ�<dz����Fؐk��
�^��������s�:�Ҟ�+0���z��d-��n�n�Ie��*e�
�K���u$m����.� �q���^7&�����#Y��I\��Z!L��u�5cL�/��]̝��<� ��wi�H}e
e��n��_��+�%!)��[� ��dٍ�SF��Gɿ�9o.�>��c$|٭!/S��]�F��*vC�JI�	�صk�VQS��*����HܸS�p�|oBߨN�P�M.����p�fj����Z����3DP��0����ʓ�w�U��#��V�����B�%�G��+*���,
οπ�O���G%�A^j�׋vb6�H�/9���k}��jna�њ)�9��./#c�5��&M\Lt���96g�QaJ
L��%�^��!8�龘ZB�g���GB�%�9�{��κ�Hբ���8ti��%A�|9=�<��>s�6�ן� 6M�ⴲD���s`�YQ�����c�^��dOk��v�i���&_�OnZ�.SrbᦹFލ�$']��Al�@!���ǡ���봜������FV�'��������0/�w��"o����ڼyϳW|M��5s8m[��ɾPen諔�(&�K;i4L4��L�,������J~���M6��i�֧����}�Y�3�dV1 o���u����]!q�� �j.Tg=���=��d��p���g���1w���?NhU�l�����ќ�L�H����ڌ4�kϡˁ&��7�B�s8�@O��ّFޯ��:� =�-���:�z�$ɼ\��d��D_���B�Ml��%�r�'{�ԣfL�
�Y���K��NHRc#�2�ˡ���0����xtm朖����H�l~�|���p���IQ�r"S���N"�A~���i���oa�8�qz���p�͌���]fZ��1��.���d��gn���)d��Xa\ߤe��&a�L��"A�փFB �[�sda{�k����uЈ q`eG��VM���FQ�Fu��C�b��Έ�VFZή�bw_����e��M�"��e�;PZ�E��j�}��+�'W�-�J��
b1�[5#oK=�,#��*������+1�jzV�G����}��O��,+�%3���fŞu�����1ov���x�x�8p�������nV>��Q7#��89����]cX?eSw}��F�/��l�er']N�\�m������r�	B�7�F��q:EW��͛�]o���06�*Rb��,��iz��=_ZG�G�ٕ���N�޹�Ĝ�I�^�5�(l�a, rK�ø.����о�FZt��j��;%��p���]�ts�27nt�,����
V����:�m��*����F�@,]7����}u�����j;�]���m׆��Ɉrl�QU�����O����o]T
6�j�49Wd6;�Q�J�?�.{�Ű�+�Sjˠ �/�/��?&j,&��W����6i�E���s�X�ŀ�9sg<����S�Ӂ�����F���/���Qc��v��R���}�����g#�8tk�$����f��8"�r@�>'<��;�u�@pC�@�^�
�K�ls�(����$������M�,T��ϰ�zϲ�ȇ��L���ƀ;b���%�g��Y���f�]��[Q�-��1�U�EQL6��(�թfU���T���\kdb��ͻ���LS(J)5�w���J���n����6M!�=��w�#Y����j����^��?�:J�a7���e0�m�H����{�R�����f��;S*���ef�����?��	���75 s�x_c�ݯ���>�G�;Oy#��|F��j�lf�{�ύ���puˉd\�lSwǋ��I�����"RF�/6�F��ps|��d��#i��H��-���DGq�����Q�JN%�L;�S����ڔ�%ǣ�+,6��:���w	��E������?R`����%�c�uĀ��+N6�4��9�T�������7�V�_5Vo>,"���2�ߘ�N�������"�SQ\��N�MV�LrG��/�Ͳ"WS䂀+���by/�T��=;��Ks��m����t�-6z���7?�e$�����/���>E_�k������5���}j@�������A߉E=�X'����j2442�I��I##����a#�<-<M���l��F���'g&�F Q������O.Pi�^�)Mut�A��޾L(_�kV���ylyF�qi���<=-�O�R�/�U)&F�����$u��x��Ɣ,����0��R�v#��CϘ���`�xJщ.��RO_��N��V 0���2��dY��Vj�ڥ��������+��j���R�ȭPYn�'d*S�.�[�R�&���=���P��ص�cOc��dP_Y����e,��93����?^�s���|>�����<�9g2_W�2CB�l8�o �]��b|�9�zŠZ;�'�hͻj/���3�~��^[ ��N��.B���Y6b��̥|�8�S���&ùd
U\�%��bE�D*�c���M?֏ B�X��)-�0���M�Ȭ��;�ڙT�J�d"7����jޯ��S]�w1�GG:���)?�2]�*��������`I@�лf���+[�<��B)���ܢ����Q�r^+j"�𷠹Xm���(��$!�+bI)������(j�k���46w�_�B��A��r�\d�q��Q?&�s �6��n��D4��Q�Ws)1��X'򤨅�+�
8t�[ӫ�SXb���������@UX'5�w0C�p�G А�ZE*F�������a]� ������^��q��p�.���	����6o��D[B�m�掉Y���k���5�z0uM���9eG��H�a��l���ޥ��j����a���'do�R?_���˾T ��韜{�OV���TM%C�(���x�ݰ6�$Ѓ�Z{��8�(�>�ܨ�Li��jP��[}�r�Pڸ���;/�,]��>Fn��
��?����_"��
H�f��?_�~*Ew�fFa�1����L�U�8���I�R=R�1@k������S�׹�?J
Lj-G�������������Z�:���FB�0� ������2TZ�փ�i���s��.KͿ.%fS��\~ig�\� �[���n�Yx��$�3��m�& ��D&C\M����f��|�)wZ;�a�Y\:/����ї��f�x�X�+�i����B����N�z��1{ �_���w�8��0�ެ�#�A�L��g����.�տ4j�oٔ1�u>��|���ɧ�e�?�kdeK	i��֪Ň���0%礴V��P��Ai�:rQ�?��hX-YC~�
Z4b�����2�)	o+(i��|��a�e0�<]��c}U�8o��\c>Wؼ ��oh�t �|�	���O)Fc3瀫�}+���,C�V���]�6pV�Tc�E2o���a�֭Y�$�t���/�l����'�ᗀ�S��ѶoX5Av�����ǒ᪷���?�\�� �F�j5���3r�!����"�#V<�\c�����X�\�gN]�V� ���s�����tpV��Ӫ�%�\շ��[N���(t쿙A,A�y�h>,֣��*4��1
�?����!$-3����xP�~a~�&΢��#����pb��q��3�N��f�����9}��<��DKA��(��]\j�����!��ak�]BL^�z ����CQ9SCg^���<�7�J�H�=��|4��,��d��� ��7�գ�Μ�y�u�J?1�`L�M��=&_F�2����\TV���Z�\Yˀ��A��j�9��9e�"8[�Y �D�M���f��`�:}Z��Wr|lq�$)���s2�φ@�n,���R�$N,sѓ�@�4e�E�??����*
|r*G_mīڇ���꒙�t��	���M���<�ɪ�f�jf��&��Cq�z,#M�0cMd0��P�%�4i���O�	�A+á���@����O�0�@����gA�}�������Z��s�a�$k�'��vJ~c���rݵ����DK�|�]v����d�� ��@���9[�"�0��S�|=�. ˑZ�pM��(szq�.�F:�\�&2��EZR�-�,���$�?H�SǀS�"�M�\��6��!�)�E��5a�L0���u��t�įP6F�
=bw�� �m0�~�-���ڧZ8���v0��w������@i��~z��se���J=Ȇ������, T_җd���Ϝ�MцCndH��#�Cm�V��)�>��dU`x&��{G���g/��E3�f3�D�$�9xڬ���F�Zm貦.O���	�b}
3�km@`��DG[�$x���#$����y�P�E�[8��Z�_�|��b���-
��`}1ZC���aH<������F3�Y�_W^<��rȚ�JK���m?��6�_%_��6��Q,w`o��l���6b�x�:�y(�G�2�q�U�l��u$����|�:Փ�Ű �(��U��$NS��+���]��N�XNX�k��9�d�a�=}���tvB%6C߰�B��0`�9lr��#-��[�b����x�(#g����=�m����k����s�/!��9 p��t'��d�7-�2�6j�!���
�#{5��ĕe����O�G?��4Aƥ޶pF�߲r�3�9�E_���@A��0c�-����(��=����oQ�ɩwJ�{+y'yAAJ�Z�Yz�~��K@�@���{fЄ=&g���3�~��Ф�\5��uk���h�G©>Y'�Ճ�=?&��)�D���.�(-�{�Y�? �2�`����k�3�q��Dӟ��|vs�gx�)|l�� } ��������-]7��,G��G܇�MY ;r�l��כhEb|;�b�\����)!��jKoZ��O?�u(9`�o���w�J{��_���La���CO�r�g���뫺9m�� ���K ���|d�ˈȴ���}����4�ǋ�vEU�FNj�U}S$9�(����Yf��v�_$Y�&����2c�׭?�/ k���:�{�K�k��S	�H��=	�8�w���B  �h����b���'M�*YK}U�B)����z̆�	4@�#Q�M \}�r�غ�]�W��!-�ӥ?9i�	\Gn���s%�X�M�}RV���6#	�)��0�X��Db�M�eΠ�*��� ��xr�����ksx�id�����K�j��;���Aw�i�=��9����^�7+��ٖț��Ҷ#����P�3��B��?_~��4X�;��k�H��D@�q �� �:�UVN �a�M�23�6IS35����ֆ���W��%���\���
�V�Y� �Z��YN���Y�!�l��쫵��D���[@�-V!��H)�J��YZ۷V-��ؐ3l��̩���V�,4�P������0�C>�Ӿ	��$`#wP=�cy���
�-��۰���澯wҦ�?9�S$����p���%jb�У�K�Z�͋����G�{�r�g#X�d!�7��$0�D���KK��]����7�,�� ��<��O]�>�p�`��.9q~e�L�+)��B��O��z�����>${�ݪ��rĦ�}�:�iZ��X5"fK��2�n�oWz^h�Ð�t�
v+��	��9C�{��Z	��	6�/����7:϶d�BGc1'�p.݄Ο�n�]�[���*?A�dx�����8�LT�@<��i����f��H_������$rIx�1��k��Vh��#�<�@��{�8��}�����(S�qp?�(ѕÒJb��}sף�F�8&��E`B>
�i�^1�K���a����S�?8���t�u2�M��"�z@�_�� j7,n�t����$�t)Rq��9";�2��[;Y#����i``��^�<g�R�2K��	�<�y
K�G�E��u��~� ��i��61u��:�v���ם�r�D��[��/l� ����b���+�'���d�n���}H��1)FTׁ��<�FQ?{��i�����g0����� y��f���pW��<�P_C,(_7�·�SY����\���	�{q�}X�
����!�kabͺ���v s�Ь. \�ՙn+�kJ����
���;1��X�vԎ��\�M�4�`?�El�wW-(:��T�?A"�m�������6�ΐ��.�{�y^��d�$m)<���bV�n�����W�t������#R�
zu����,��,���1ޕu0��l[@d4=�h����z���P�i��e)���;G��at��^[m��cW�kq��mZ^蝄�<b��t����\4�G�y�Z��b������*uy[�Y��?K�DS"���P�eM��>.��oV�Ꙁ+�H��i*��@��ϔ=��B�q��<��I�v֗��:g-��y*���U[k>�.�V��̑�]��U{X�> ϱw�.~��ŗ�2����E�.N��Jv\���(��5mn�T?	��b`�&D P����Ta�Ȕ��^��Z8DՂ����^��ΡT����:3LxG��g���Y�~SB�P
��p1��w�sL���i��5�> ����J��/QM}������Mln�-������o��b��D���������Җۄ���J1�91�&/�S
�Y�·[;���j+����C���t�cz� S���.�����Q�%|�z�@WV��~C�œ��!NC��0�GY!�C^��_K�a�]�� ��*��J�3�R)>=�,>�s��a��6��f��ne��0G��(�^� Xc3��Hb=��Nd?��+��"�Z��Sr2���ć�q,xB�!���38�.�R-I�-(���g��4_*R���S�����Ю[��=K$p���eBa�)7�\(n���o�i���hi^�ILN�)@>��z��~k�2�����U/B�4�@.�'��˖8��$]���� �PIt���V�9���~������NΊ�LU��I[*�SN�K��N�C �j��N h#f�FL�Edi9���ޥ
˨:�@��ҭ�j�fj�S���B.����6��ץul������b��76x��r��P~.zL���A+ٛ���/e�_�U�綱p����\9V�Ҝ���4�m'\�%u����'���!o/j\����ÿoy���^My��G_d8h;�o���-���"ʚ8����'�&T�&�MI��9��`�ޡ�%ʸт�S��>��bE��;�C>����1�d2V�=.|4�-f�\� &�xʕ$��D�N|�����*�zj��?l`�~�Z��EȜi�/�� '^�;H��Eќ��/�UZ���7S�S�����{�ظh���Q�����˫1��}���K\��?�,�:*eM��!-R�%�nW2[�!���������B��T�yl� -��e�-��m��瑚Ѷ�UCh�
�3&�Cv~W�E_���ު񱓸��cp��.É�� �b��r�}�,�V�7�~WYխNei�]��ӣ:�lI&�X�J������ǵmЇ��;A��<�.��Q����Yd�:�
�%3��m@�yCغ7��㧱��2��lCC���R`V�w����BB�9�􀇗χ�`���՞�g=��kxn}᪤|t�Y����dAvI���g�ݮ�*h��
�7�>X$�3ະ8P��vi��(�LK�����ھ���W\F8��p�Np#��AwC��sĴ��j����q�I�E��:z�>����FHb�n�GS��y�E�R�t�J����O���Zb����p�Y ��o�7՟���yr�p 8�)�p�$��3���N�a�~z?����K�-��������x�w��V������񌚼�.����f����PK�X* ��0jwA��b��
M�C�J������3ป�*.�Y0oY@�u�٠�4��$X���G'��Y{(⋢:p��3%�^��Nf�v�z�P��A��"�l'lE�;��Jē��|s)��\��9n���_f^$zs�G,߽d�hR�9$�3��Ch���-���-�����gb�a�K�eee���d��ץd`��[�I;��`� �}O� ��HFx{f��\�\-'���k�佷�x��0^�#�ֆB�vtt\���v�x�4�W���F\���j���k"HST�	���\M$���~��vq�+%w?[a��d��%V9w(m;B��/�Q9D���YfU$yi�eX���hP$è����ג⊊�fX$��V:Û򂮜����<P�
�,G�/`q	|�̟��~X�,�JL��rA��چ������J|b
m��H�e���t ��K���?��6��~�K���3�@+)��f��%��G�C{�A���$sd�]f�%]JJ�R�SOi��q�ȇq�!��qP�i�_���ȼ��h���88���-28��z�6b���+�XB �ўJ��͒>�w1��e����q� 7�wZ�e��)P+STTb�����Ҕ� ��.쬝΢0�߈qUڝ�2r ���Ӏ�]��@	�l��\��~�,��k�M�;7db�kZZZػҟ�.Nld+�3r �Y�_�R��>� ��ޗҳ>i���V��Va�1D�E0�kϭ��a�����EC� 4���DE�A#奂v�J�a�ڤ�U�3����x�К"���rに�srk͈����y�P�aH}k3π��S��
���{E'��t��_C�Q�g]9�\J`��G�ť��lL����r%,�9U�����͏����U�M�]��#�1܆ϓ�8���6�:�FM���@�Ȧ��K���>��7,��?Ö�,�1��[OU+VN�)?�$p.�q,��U������P�����,�9�������:��E)�N[��=�K�|��C��uL#,�����z�f� ]�PФI�0�']�ʹ�e�g��z=;�ٸ��Z QhB/i���<{����������hd��0����9�����*辪�j�ӏ�|1���Ɗ��T��� �k�Mi�z9]K��}πG�RR7�	�㭹����ˮC3��άUY�%� ��)���;ef]b�?���2	�����6A�����>*%+�֍�j|�y��Hܣ>)�3�Pf%��JSo�~T� <�=W���j,`�Q��� "E��(˅8�`bb��3޶w��J�6���c`��^?^�);qV`]�;���M�p"�� ��[��@���ʡ!{~�;	�:�/l�{䇟�[�Z���Es=_���{�=�րᯏ�zP?�SA��d�*�>��"[�7�^��%=�<D���k�������"� �[��%�Ƭb[�,�7��U~s
�P2K9[}V�wƛ���+�6�M���+2�|��M�ڵoƊ��4K����IY��X�P�|���Cc|m\��2��5Rzn<1�/:_�(A�AN����K5�r���z�#e��b���\Ȉ�]�fK����a)ω�iLi�Iݦ�Ȩ����Y����n��4?��U�5d���N�W��UĞ��&'�p�+��D�GC� ��q
i�%F���ٰ�z6�'���B5�Ĺ5��W�3԰�,h�w��e�c~'�����"_1��.�'�����	�
�^к��c��d����OQ)Y��sb"��7�Ŏ7���Sn� $���e�yVh���IÔL�����(8l,w��X�ΗF��u
���q@NG�w!�g����l�z��^O�3�{c�<�N}�e!�U"�nZ� �giK��1Il:o��3K���Ok�=C�آ~¼ҾT�8f�:�M�(z�mL�� ��bJ$�$u�`��M���Q�g�k���2�g[��6�ǥ�2��p��[���%&����w~�B{=�&-��N��f���Y�m��s��$a������x]����(z	_���jϙ�:����BM��-n�I��#�G�`�6�z ��f��؜������(��.��1 ���Ng䅣�3G�D��A���'1��Ǔ�'���
iU�YJO@Z�נ�*��,�X.�MR����=6�f/o]P���8K,;�����H���=87ϓ�48��d3�
�\Z��V�E��<���Ѡ.����5SWF�՛�ڋ���oa6ܨ������ނ�ٮ�M���?E��Oʭ��0{o��:A(�O�*[���7_��,X��DȧB�w`H�K�R7ΰ�����m�f�ΐFjir_h��w��.�����=���TjZ���%�)�)١�����kJ]|=v$�"�t�.�B���(�d6�q�ɦ�0�'_��[�X�����k	��S1��n}W�X�֐���>��ڑ�W6��K!H�x�N��|��̰�jf����q�C�`����w8vSQ1]��+J4����:�^� @B��xX�>�O��8,B
89�nS;i���k8V~���[P�GGG�0��Č��a�E�<b=h�$���>E1$�%[��s�S�v���}q�5��܈�J�R�ܐ���$��e"H�-Ѵ�5�!�~����*}~��F��(9RӔ%���!��.�VT)`��_�V�����/I�7�b��a@�;o�?V���<���������l�Ѥm�1&�~`idd$�*iP&�E�cAJ�����U�<����� �`��tZ���z�U�8�Ջ^����/�=�	<˩x��T3 ��N�k���G�^�_kB{z�h�FD ����~��,���A[̈́s��J죀YX�pa�Z���U���d�N-l½a݆���7$�B��'v$����x�!��Hn�If>���Xgs��%o}��"p� �,2=5��s���s�%�)�#�rW��Q�����z��)�b�Y��>x>Z)��7G�y{F�ft��złA���BP2bޒY���& ����@���$Y��r�	���V|��F�n%��B��t��$@#��#-���0���v�?=��c*q7S��=��qR���O ��n�X��ϮZ
 8/���j�k�`��!���Ub�:�ښ��TOϜ��+���SF�.���.�a��(H���+�~�9M�7�Y�BMRRU3�Dce�>�RRcaշ/��봣����N�r4,���D���><�l#��9�Ÿ�]�4���T˘����
y{��T��>���/Q]���F�-B.B�NSKl�DP��`C� �ч@l��ǳGǹ��}��齾3zL����{��>E�}q�,53��y"���3\=���������x�A�}c��?�k{�s�ob�f����
'�#�%���b��7㑟�^>!��PS�j4|^d���Ic�J�@�x�L�����<�0���j�Q��5��^`H�MQ&��4�!����O���"�ow��4���q�e��m=�aV���W��$z��<�.&�UJ"iOVti�/�����8?�1�2�4�j�jW[��lDr�䀈`�1�/���&9%3IX�
簫�X��i�Y�qx��G����.�y`��g�{S�e�
Jr�5�>�#�җ�NƜ��2���'�
�(�u�;d�~����m�ˌ�b�	]}�!� ��t�ϗ9�9�gv28���Jf�r�����c�O���}u蠗t��!3^KH�os0?��*���Z���H�&=9tUFx��mUxj����j��j����kϮ¬����>�)@����Ƅ�s&+XL]�K��Ģ�\ϒ�F�ӏB
@�bN��Y�#e�pR��I'(��fr	ܛ�K��[yثT����d��}�lِ�O�x����3��;����888(�q���^�5��(*Z{�.Q��L��v�������F��@N؁f���\�%�|*v.���rD}�PɌfPH�{�Z�+��,��і�>���Ȱ�mmmOa�3�ᦑ����IGE,8�B�a��c&�ډՂ�:�\�H.�{F��%l�K\O�+���d��ؓ�Q�T�q���SlI����A�!ۤ�u,�"�˓Wr�;�a�^�,H��M�U(��ݰ��:�����F7>���&��ʿ@��L9
j;vBK����͢�cW�|��	���{�_�y��̜=pc��� �8���8o����%�`�f��{�����a܌�T�P�&�u?{����cb];�	�J,�X�����$��	��iry��.+*)�Sҽ�֠Rŉ���DX�7��pQ�J��$(a�-�r�>Q9�o�K��o�����BAk͵�� ���9��~Mj��R�D�S�4����ˬ����G��R��6)� ���5�����ƛ3����`<�V�u<3i,�ڵ�"خ�.�
��-��>W�ڤ�6ň&G�M	�g�M?�C~�U/I����Gy"웽۔i�;��wן�L���Tg+��A������UMu������f/�dH䣝��~�lE�9����d������I��ڧ�N�*�|�;[=c!J��x���	E'*PG��U�}���C%������k�%���j�)#e�SUS�x���y��Cu��'� . �0��;�fĥt���Z|����oR�mU��C��7"H��
X�exݞئ�J7��H����}G�᳣��a>�h��WD���i�@�����@�ދ�	x����kg2c�n���6�q���
z�������n���5?�wǙ�ҍX���W��V)��z�՘
,
���%�U��:���`fcס�l9a�j�5T`?
�W��+R�%�K �N��(]Wr�*W�]�Ӳ�<7�E�Ԝ������ �)�		eNa?�h����M6G��k}� ��n��pn�u��x:-o��ްc���B�d�Uw/�`�'�>#H��Wb�sJT穽sssE111j]���l���ۤղP�'}��������4`�,��{߬7���+m�<u�1��T��q���VH�?jP�̯�;z@�%E~f �V�+-��G���^�zT8��Drf�O��sF���'�D�Ϡ�߻<�}Ɨ&t5��x�I:Y�/�^綆>2�8�;4�i��ſ{����P͝l�\�(�˅�/%�� �
pA<�����p���&j�x��˫�!��&J�q���.o��.t,]Xdu�?�w�*h��Q�[�����3[�N���a��w�w�sm���ܴH�k���4fc����9��Їq��1�S׀㚺��|� s��\BdK<_I̟��F?��r8u?8@.��]]�3����
ٌf��<���ޘ
�k����,�߼�ؙ�}[�e�G��ӗ���B�h��!ޛ���eH���;~R�9�%#A��|[�&q,j�~yр���w�|J�� ��������2
��bJ�u��;���>��=?�{	�oW����
������^�o���G����08K4}M|���UPo �J�נ!cA��g׺Oչ�h��-��|���B�Qܓ�ځ���i������vx��m��I���*f|��D?1W~�W@5�vdr(jW1�E�=�k��s71�` ���D��D�|E��P��d����Q�$�j)�+ӗ�?ÚN>�:�,��H�<��v�w��.N,�H������Z��V�
yNOѽ�z��S�Ntc��x0@<H�J&%wYsEtf2��ۅ����dK�
)!^W�����	^�PF;�?�׳U=���m؏g��v�5�w�|A�����1d�*R_U����<�c8;�vCl�ގ�\�����o�H,M�`ŭH ��RF����:�N�!8reen����;sd/.���a�J�v%��� �w`,>�e�����y�Z�����@�G����N�H�2��Gy�(�
�!��Eu���e���3��0�.@SR���@������Fg��N*���$���}HO%|��W�NʜQc�� )����Ǐ�V�HZ�#�QO�1I��A�� M�M�O*�Y6��?VH��G�Jb� Z_�(J��'����n��G
[� 3/�j����;+	!�
[��B֟�:�%�}U��
�l3�f�*�(�|x�̋�Ê�y^A���'��P�?!�xy�(߁#}ԅ�2-D��c�X����$�>��r!��~ N�҇O�C@x�C�xͿ�g<ƀ�2K�x>�骽�(Yܹ�>��gb�^Y���0Ot6eWm�gس��u��잛\J��@M�1���
�M��д��*.�Uz�@�;Н��ff��pZw26�g�7���[��1�SR���j|B&������/��p"��*������//�g���x�K�+*sK�b{�y8NI)F����W�7��c�v��� н*�u�����r/`tw��;(2���hVkԩ|m��>�?��>E-��<�> �F�Qi�|�
v@�w���P6%2�B����;Mps���N�h���%Ǭ��r�ĆX<�#����\:�𽦀����='�ۄ��~0>E�Ja.�D�W���7��J8������G޲=@�wZjs���N_E�!bC^p��<�5J�L&S�{ei{@H�	�"�*��٫,�KX����h��Ő��̰_�M�Gu��>��1�)��NQ<PNޠ�c�"��y�xuwbt�UP3�ٔ\ӟ	�u C���0�ί[��i�����Rk���Z{�4������G��J��w�~:�f�����%.N$a����l���B$_�,�	XF��	Y�R`����(�� Wq���_�ʡ�K7!��N!����Sv�O�H�]�%,����`�&�xx�����F�B�(Ȅ4)���~��f�A˿Ïa��5ԷCP�S��2P�2`�Yj� ����G��j"�jR�|�ry)�\�"àEA*�,��
�} �����*S �*o�bO��� ��c����\[�߇!ͰS>�,�J�����W��Id�i��u^GH
^��?���$�m����4�՘�斸��N��k���!�5�m��'��81���Q?>4$��p�`��:��6�*!l}7�Qz��t����R����8��9�Y�P[�o�[Y9&I끯g�F�ID�_�SO w7͘������%�p\��!n�=>)���M�L��%�� >����C�����������Ѡ�������(��_��R@��3��r#;FC�gi�#
��P���o�}�j��"R%ol=�Qi��H!<&0ï������I..�h�CH )�֛��c�r��CJ=�luM.	��D�C�l�OL���,����Qw `P�.�ߧ�\v�5?��j?`����E�@�~���O~�ɲ�v4߽��֜eӆI�c��9,�A�7�G�������ܐ���S�Г8���OcE���ܹ��>� #������FA�� �QT���!g�D/h��Z�%�|6�9��6ZYA����K�����X5^���s�>���E׆�C�ۻ�A5�{�m�M:�W^R<:����8�����hE%dz&�%=��B���v2u3�i�TGa�9t"�;��4�L
��4V^�mA=d��п>�cA9t���N���2)��&�|L���y�.T��il[�����t�G1|�����5,]���s��x��b�!�sӻY�Dg��O�!d��E���!��o�烾vJ؆~��f���6ĝ:w�'�n���!����N��@^iL�&���UYޮ�E�/�*΢�ubo��n��Q���H�fd�t2!�8��������4L�.�V�xR����YEI�B.��8��C~3`�̾����R���RD��0�E�sֳ����y�Ri��Xj�mwOO����J�gC�@�؇��}�������i��_������f�׾~£�a����(����q3	� �z�1�l��J;x՞"{�o?1Qv�w�����	�+��8rs�n��+���5Un���M7!k���!<^���ċ��V�t1���,��YB9t�%>�D<|"OPG��s4Z(�PNC�PZ�;1��k��bib�߾�%�f2�����UI����Z[ZZ�:\� �:��4qK�V�-9RZ ��&,�;wN�|�����{�*�bBi�ӳ�=vt.��Sn�Jn_��F���M3N�1��
쏅=�T�����g�������v��u��Z�J�9%�p���	$�c���\������;|o����F���jY[[��?�^���fjb�pʫ*�{E���o��옷g����Y�'���O�.����}��0� �8�t����ɬ�X17��&��Q�,���R((�ɑ����O��eeKx$?4	�W���E;��{��pM��xm?�\����:��>�we܌�*�x��VVO��T0�	8y���\qbbbe.�o�> >��
��I'�;|�[�$�X0ϩ��k��z\JX(�ap�D���M�[��V��jqtҭ�oC��]K����������j��R��D%�4�À�sp`�א�7��\d�]SWw��j�%+�ؕ�q/Y0O	A�HP������OԷǥ���I�Hz�%��5�h���*~L�=�!�,�A��}�;~U���W�?m�
�����)�@��x_ �?=�-!E����'!6JY^A2�	���dX�R��!$��nD�O����a���}��0����ƃf�@Sj��x0Qk}5�QB��%j3kN1�R^\}�"�I�p`�� �*�@\��'���_��-)ᩘKo��$4` ; @&p���.�z��(��@���{���-�7�j���+:���ÇUٽpڜ�M�֜��`�N�-�j���d�Pj8� ��`�/��a̯�&�������fC"���J(w����������*y-����d�'�}y����@}��������7��ڡB���X��'*jI!80h���9�3�l���*��?@���K��*�q>~��0]�ꓭO�w	��΄7J�7<?���eO;����@��)Vu��m߫�[@����NS��U��;�4���%��.9%nO��)��&O2>����j�_�� ��]>�ܕ�M��T�q1����
�$�V �&�Ŝݞ����_<�;�;�)����jN+���M��7z���.N��V~P��哛Vs� %g�#J\���IpI�2�;�֎t��Z��-v;��}	>s��l�nHopXs�_�#�/�~)�����,or�'����m8鋟Y�i�����������y�ж��{�5��?�Nw�Q����-���h�v�p�_�Q��@�M��c��?��Pt+��\��������c�
�/i)ߍ���٥;�&������SJ/�MR�t	�7�WV����s��:��+pf���K��.�8_������|lg0�m����к�_-�7|�R�&�:�ۖ^+�TmSK=���H~��������\\�n+�Y���ĕ}LL;��S�t���]����L1���&V�hM`y�oʙQ�Wb�>˿�Nr��PcS�) ���]�)��s>�&.D���	�����i�.�Ja�4xݸ�Z�۷��o�O������ŷ��ʦܮG�>��0*�U�^g��a��n�:t�6(xk؁b�*�p��z��%��`�2��B���u-}��ZnzyW���O�5o����~��H*���N�s[��C��	
�ޝ�^�뵁���|��p��R������y��Z��o��w4&:z��䭖4�f�<hʣ�'�ݼW��[Fz�餯I����'�!=uHW��[I�c�g�mBI-����b&�/o�4����r�w%�q���w3����t�[`�⎬n��%�VH��N��J�{Y���O��6VD�(@z\���b�f��ү��o��K����@�F�����y8aSgI������R|��)�`�s��G���8�yr��y�9'��t�6���N�Mu^ʅ��;;�k�TYBm����vu���/V�oQ�D"�V��<�P2��4q����io���/-����þ�9���v��w��yn�̬�T�s4K�s���|]g��j��Э�;'�w�0�<Vz��)H7h���/��35��j�de�ZU�/�v8�o�w{$4b%/��i�;ׂyYd��+G:��y��碯��|#}�%�G`���w�v���<V2N���2����Mccc�U.�HV�W�k߱���{��T}�gaч��Q�kd쳯��K�-�����}�RK1�"����XA�D��q������N����|�tb��ܴW������9
�yTn�X���J�q��
k��@�?�pN����;l�h0�M�V��uv'�hQY�>�?�X��iz��%��?m}Bm���}"iT�����\��Y���2��Ƌ�'X������{1�Ҭ��fh��*�y��%�^XYYI}��G4���AX�랿�k;�Z�5޴ggx텈���r:�g�%�1-�e�r+��ǥ����h]xF*�]�4<�.+''�^�������ź�+�������L�W�K����+ߜ������>K�^+���h]���Ja �rr����<-sAeȁ�r���*m��XX�8���}n��%�F9`��c]�l����9�>�3���d2��VV��m� ����׾�nv���o^�M$�0��ٽ�r�L��Y����� �(�Fɱ9��	�륍�����5�=H%E��$ge�|�k��?�; doǏ�1����{�,��ݹs����>n���l5��󵶳��Sͪ����/�)?��>`y)�2~6�{��/�|V"_$��A�r׎)��P��am�yQ�7ͺjTq�䗄�A�w%���@��f��S��!=�N���B-�om�6n~&��Qf��k�w���;�Vs�� ��k����n���@���ҡ|R��o��{����_��]]������E�M�qi}���cx�]}�q[��� ���t��o��쾛���M �\��v�����`dd��������[䵛{}d�o�w���k��Φ�@��]�\c;�>�(TZu�]�j�O{���B�fE���M��7�#^��>�X�qǍNM9�z��������g�o��J�o,H�< w�색�j�b�B�%��P|Kw�gC���B�����	�RI�a�#�<_n���<���"��I�F���\\!�����5]�!�f�|nTh[���-96�Na��nUUT4�v��I�l���p���L%�l�����o�H�i�R�p;��oGt����F��v��wX �[z��'�_z�����)�G`��P?��i�X�x�j��v�f��U̥ٽ����uY�rRT@����V��\,]�t�]�qO�Y\Z(����n49��x�>/�7��y��0E�z�ݟ�?�-��0�~��]x����)@�q�Ϯ���vT8�]W����,�$�84���㲒�^y�h�6kI�ke�p�;o���#���a�4���k�Q�ht�����eSDˆ.����x��G��&�u��B7�P{��,&�[�B���0xpCCdܠ��B��w���#�ϥ�Hy4ix����Z�<옱��?�ˤj@A��GU�@��mHgxvtekG,�^Z�J����DO���׽��`�^F/�$^�T���A�۷�b�M��P5�ɰ���.������
�'�2~�Q<g�b���j�j��]��mz��|�KL7��0��Iކ�
oo<>7�X rɻ=I���{>��W��M���a����T�x��5����j��c0��ݝh $7z������_�-h~l���$];JU��q���6��"d�߁�;ݸ��}t���ڏ02�����O}Q��/���kl'%�;2�1��.F�w!���)��4�`���{aӞ����~�xg�.����`A��ۧ����:lJU��"����B-Л�k�p8�䉮=��ɋD��+r�x.���o���S�\��=���>G�Z��?���@�T�MP��;��]�m�?h�73H�~|����Ŷ�J���Ax�R����N;���7� ��_����r���c��zdjjb�<���a�X�Z�v���I)��{k��e�A#��3!&�
b�l���(���;R@@�`~����9�R �M���J�wנ�
�2�:���:?�N��%�S_�u��9|����U}�����>JL$v��4}��A��c��j�~}c��Yug�ȁ
0�~͵Ϧ�3��_�
cFGh��d�=<<*F�&����휦|�Q��e�[E��ϴ�Z.�*xʼw�����<�s�״�}V:^�D��s�I��'����`�"h-fp��{��c\��O4P���eL���D]�M�*��NM;����]>p����HOʣ~1��nĉ��W���]�J� �@��~�T��7�&P�?��E��͕)ߘ�y�V���A�c�r��#���U'�\CAѮ�^c������Ai��{����@����*@��_� �m��nRD�î�6IZWIX�yE��s�b�Z[U����@O��T�C`R.� � #�|�F�BDg��c���EGs��� ����������~P�&{{{#1�9�@�x�|wbk�m>iӞa��"ݠ)�r%���I�a���-X���4��;�Oϛ��͸�-�8a��3D����|���Lk��X��R։����\MMM?&��$eBr��$][���3bo����d�_-//�z�f�-��ǻ�{���e��K)���|�"\�H���\���5<��� )7n1>�ip��Ӷ�e�1
0��,�䭥����=���ǺUz����D4�v⻤ݜ�Z�	�B=��ȱ�1ء��i)=���(�0��UC�U��C�3���k�����56�"��*s:��+����m�`���EwF�����Ǘg�+W0t�h���E�=��C)����7�N�5>ǧREs��,;4~I��O�TI1y���tM�~����e���G�����%�T�m��P�H2�
�� T2mlIi24)2�d�2l��D���XGE		�mI�2��L�6Ŧ��?k��������w��:�w=�}�ϻ޵��^-BZR�A�LTD�mS;zyМ&,_�)L )�bHQD��I�;�Z�L�
��I�o�ԓ#��}��d�3�([8Jg|Qa~)���3��S��Ī�L&�vtx�b� ��t�D�/��́P|�G\��J�l:\9��>��߫��BJ򗩊_hƋ�����zf�<�P~�5x9��I&�`�#`W.x��,��8?��l�A����լ�p�;-j����u�6i�&n*��O�lL���m'o�)r�L�� �Mc���t�=�=[�t���M�'� �H�ڻ]�ˉ�������֕��$�h_����Ҩ��e�tF1,xc"�E#wH��B͵���i��3	�$�!w�+� ��
;5����o@�S���7㷼�͆G�w�%}y'��ۻr�@�^|��c�k�`���f>���餜����pP�Vvgs�
F������}�V��~�]�p��Z��X�2��/�e�uZT���q39��l�� #.	�'Źԟ>O��?�����hu��)�d��W��������z:\�nͲ�E�x�I$p�dWy��ŀ7�:���]���ng�B�o���=g��^�|Z������=�+7	Ġ���-���IH�����݌��ȓ���ӫ�e�
h5���I�ze�b�u�t����;�����ga��Y�H�����\�*�I�)��_�J�&}U�U=Z���IA���� ��q)"%��5�t��a5t�z���0�F$C��|8����Sy�-�o��*~�A� Ì���N�0t����E���~�Rė/C"�;�8�m�<�-5�vi��y�}��+U�K��3��a\�FkS>����~uA�`���˗��Xw�t��Uw��/���{Q�C�5\�k��Z�+g���&��O=������e1z!s���/������r��S��S��yk�l~ߌ���d��v�-�l��0���,;4��u�O�r{����h۳q
]Gw�����`F�V#/%�4_��!䜢���E&���dݦ�C;As�]$}wtt\�~��}�լ�:P�oϨ����U�y'���w��&�b ��.�1K	r|mQ��
������|�÷!����޾B$}�D�@k[��Н[̞�K�����*9��l��q�n�N�n�iL9�W��˅D���p���C�6�3�Y�OMg��t���5^�|7\\�AO��ݻW�-��jˉ5��_�.���f������u��,����w�x�*�̷fQ&J&K����J��	1�O��WO{s�pn�g����Iߔ5^��M���y:44������m|��c�u&'��Y:�A_����aV�x���i�����ȏ�#�*�m���wOVF��Fۖ����L���;���y;3�+,:�]�5���a����gO"����R��S�\�K��*^ tv"/7�\TL��J� Z�AR*����?n��D�teGU��ג�@�[�P*#�����5�Զ��ȓK��-yj�C�K�J(��	}�����B�����g&��q�NTWx_���pi[$3/���H�̩]WJ�u��?3��Z7��`�Q��3�EPy�x=s;����l���Ձ]J�Y/٩.���K��a�����]!�F
G}(��X���H��7��ţ�GM�VT�|s��ן?c��@�<#n�'������79��=�[I�LLLnCR�>-Ss.�����M�:p-YqH�Q`��v
�8�b�c�]�JMA�&�쒗��ҮO����p�V{G�b��-[����}��9|b~��#�r22���>p�U����H_�@����MW=�z��,�hZ�kr�+��n\��u�O�8��T*�MV��j?�� �+��)��*vsf����r扬hW����-ggix�s탉B9#�{�i��o|��1���-��LS0d��S� ��|��M���)>>~�g1٨�3�:�E�i>�E?=N�x��?4f�͈��㋓�9lV�G�5�P�~��3���E���_��v����šai���1�1}���P��>ע�-}�4w���R}���L�o��(/�S�����|�~�&����3TS �7Z6�@��()*�m��Oݽrѯ���ԣ�����C&�Ĭ_��*�����/�yzz�N�4C/�7�;b]���^_���l�B>qo��;m���De�w:pv?�Ӣ��[b)�y�oHz?��J���=/�V�W�:ǰıv���5Ԗ�C��a"]���Oވ��Q���{�W����w�fR����xs������b3#I�S˹��r	��F��Y�N��j���h�������gB��eGrֈD722Z,@��~�d�jt*���͑LVB��3�b�Ƃ�;�V��� �;�>���)[�;)�XL��o�Ee힡=��[a�V]�%���|��� /���,(��a���_󅃓�J�S>}�+m/����π��k�G_�e6��:�;}>���F��j��s���G)GYi��N#&6
>��{�<"8Į����15���>Y�WTW�%tQ����﴿oM2�-G}�_�Ʃ)��a:ݯL�%2�k{�7����8�����E����dQXg�K�W05��[c�w���S�^��91z">�/j��}��c}�*�������h\/�����>�i�.C��[f�P٩=��?�Jk
�	z]|r!�^I5.W���Z�k�=xBӱy���Ƃ����'R�������>��\��*piJ=,��1qL�o>͈d\�59�G���/SG��p���E�����RT��-��Ȯ��h�?毠h�<��eA��@f��#�����H��%ޢ&8ufo�ay=���%R� HJ��֧�"1���s�(Z�Ow�m�;�{���c)�>N�EGb�?*M�U����1�������+�sWxcb�&������	sƿ��:�m�V&rؐ(��vi��%G�����*�_���¯��&��Cg�>t5�D�R��;;/Cyeg���|�y��S[I3��}�7�Jک!Q�$�X�d�yi{�-�t�M$���+8�!�8�͎N���9��(&��<�k>��,'/oι��*�������䳝����:~Tj�q���<�cv�(2,QϚ�4�5X��M�wJ$Q���M�ԟ1av	'w0l97�æ��Q�~:S����M�+kn���ʧ�R��.���݀�C������ː݉9���0������B�w�[��c���N�_�I~�G'+�l��\��x�r�Ʋ��q�7��{���v�'<�bD��Au;-d�X�n�����7hv	��|_�DI��!F�*�m���T�g9�Q��/�fH ���\Ԩ�m��?����)�-�RW��(���fF}��%ٮH.�&ek�,rg�Of�Nwб�����m��}xC�gH��CR�i��:Y�f,�#�g�'m9��}�^�^P?�=�y*A0K?�5uys`N��
+����jj�0*~���z�Qޓ/�S5np%�ŋ�wJc���q��΁��:��.�ɭ���ԓ��I��!��n��'��ɯ����e�#�?�hs�M�i	����i|�����7o�ddd����@��u(Kڡ�Evj��Ǻ��m
��v��U���tΑs~h/h!�R�:S:5���;�q(����yn�J)Q������s>D��h��X⏬p~2ğg~�|�Ľ��:��i�||x[GGJ4v��d�|u�'���W�1o��xo���FS��ʬ�,�Ƶ���Ԓؓ7����n~���#���i���R=>�z�q���ki�H�������&��boRu�t�+�Ή�&�Y�{e?�m�*P��e����g�T�-�͛�X�L�G �%�;��4�U��].ڙ��YqyiQUs����ii���R��#AKa�X�m`M�$��럾�1<�l���~�ț��Ҁ�@�侕�G����Bl)�]�����-ڋEńɲMؽ:���n0J������S�7��z�%بp�GO�۵�+�%n�?Lic_t�Y��N�$�'l&72�.WǾ�N��K����zdK98b��7�M����t:A1ث�����'��]���B���#��v�W�p��ˇ���t���5Je's쵼���Uu)�\���!�S�D�i� ;O���$��7^T�j�4g���ϼ_��>C��30�6U7D�˾K[��Ȧ�i���1��*�6^��#���4L-���kl=J%�9�  �4>�Hr�R����_���H����Ew���~��	���O������w!:'��"���L�,���U��ɒ��K �$_W�?A�5A�Y�#W�(����$�S<��M�XT�� *���5�.�8�r,�$�p���(�K^9����WA~++Z2��B���tG�+ڻ�9ө��锫#aW����PS/UZ.�,�h���V������OU���Ay�	�P�m�&D��=%�uuw/E�Wt.[�d;,Z��b��9D�y�������V�=T�m�ŋ�[q0\(iJ*y��D���P�E�f��8_���b�vb#kv�v
�xbfױɭ�j�����B��NY��,�$ߠ�^{�]���	�U}�(���>���C^^ L��x��{M�%��ɑJ3��e%���������x}Z���0�O����d�Sbs�DJ_تʮ<YZJ�@I�ݚ�A���^�L�R�M����E~H�W�
�V4���=�	�I���jI��6�_N�_�=M�'�+��:���̣X	U�����
[ZZ��)���½����� ���
���p��Š�d
��r��u`+�M�-YDGM��[TI��ꢷ�0��{�h	+E�/��3�%&&������Dl�K�4�7�q~��̓%� x��P��4�Ou�b�.�
��R���G�<����cK�=�.\�&�>&@ƴ��e�c�za���U۸��aZ��p�@KFu\�vB���3_�׸�ǹ���^���_"����RN ����·���$Z'yˁ4a�����1޶�C�mBgp9�^������p��҄�p�'��+�/_&�X=I�Eos�t�v�%��
Um*
�𱾾�<N�w�ce�ؙ,�}n:����3꾙���P����>��\�U�-��o/ٽ��[q�a�!��<iQKj���#ݽ�G=XLt9%x��$5�ϭ�e��Mid���B������p�,��Q�2y�.Z���K�;!�傴�s�v�=��t\\�J"L��BVJ��N<6�꧀�ɲ�DP�
OTvqy���U�.�?g����7��fCm	��Y	���O��+S������2xD�w���Ic�=��_�\8,���԰Sk��.N�u`��5�[f��,o��Ud�f�Z��I	� �g�2ݙ��3���]�-�4�gw��u=��]k,f����&���n'�	��� s�K���8u�su�B���#����CCC4r���>0J���c9;=9n$��)X���V���hO��=2�"γ֙�޾Ђ���''��M�C� d��xkb�}�,ࠇ"�P��;��=?m�f 6r��MX�J�DlK��֭[y���{o��'ҰV��vn$�]��B#��(�6 sL�^V9��~�������f_1Ά��H�h�{T�_H���o��� �]�܀z�r�����n!���gJX��Ӛ���o)x3��B�e��E�!m�m��4ՁoC��ˊ�(+���@yE�'��ow��=<e��t����ȵ����t�+\��_<k�M`�x���c0lx4�������	`��=ǿ�����`�y��E�������e*2,|�B)��8��p��a�H�雼>����P�%a��]���J��o���ydX��RW���̍��A�����ν��F1�x7<hL	F�Rz���i�:�p��ҹ�9�pt�x�r�0rq�G�\�#,�,��۫�6��I��n/�z�C�da�;M���-�mSCF�5�N�M
���ےdj>�(/M����c�m��D2�@{�!���[��n����;��2P��T����?;��	�|�ˏ-�U�/�4q�t�S�c�ɧ9��-H��u��Ҽ���Gg�u�ۼB�đGU�<�GV���%����Q�n�By��+�,�,��
Q=���>ӕ��y@����s��^����OU��na�V�~�E�Uʖ}�T�UTL��<�Fn�`6��;hοG�|�à��.���1'`حr�~��߄X�Hĩ��n�M��z:+�7/T��6��q�a�{��#)��DU�AP6 u�.qJ0δf?f=��{EQ�2,v�un�,����������x<ӿd��!��c?&F�7�z�*,U�n`W����vѯ�}��"g7���y��,�����~�MbqQ�����F^�;m� ��������VC�F1�����xE��U{A�D�mh�t]�����V�������0�@TΡÙEX}�mY�J�cX�XA��(f�<$���{�gBdIKޠ%³Xȸ��e`����q�N#��ڎN�PWaV'�c��j�Dӯ
�3�;U�W��66@Ex������z��`��*������`H��%���uV��Ug,�:���~���!B$���e��E7��NN�F�� KX�O5��mG70�j[��4��d��A��F*�t�~�h��޳׉��|t�tl�m���^|�XL��:,fZ��\������6c
J�(�ՙ�x����d�B�ϴ��/9}��DAц�aJiQ?�㭞\�A��{�z(R��<E�ր���"���H>��u||<�����@���D�@w���ė���;:�`��DrQ>����_�����ax�"{X��t��!OW�>�%$���/�+7� ��u�sh�����2LQ ;Q.��o�th!�\�$��yE_ۍ���M'tx+���rh�z���)�M��F1�D@���6�k�f]bIAA�r:)�iT*��7P�����X�wߩ��-�|��P3T�r);u^��~SnQ8[Z�����]lq[H��<����<I��%����*Y��^AUxҗ�'�F��R҈���8��&���7�ܼ��7�%�]�:`�����b~DЅ����E�� Pp1z�[�].7�g��#�����l`���i���.)�l��<MJ���ćXg��������[�C��Y*AA����[����}�,i�Z���{�y��ԗ$L����,��h �6	�(�=|iȥ�F Ф�	�HA�~Ɍ�q��eґ�*u��~�����G���'��UB�>�;�Y	��B߄7��a�wSL����ms@�	<�<�<��-%�a����|J��(�5S��X�����hC�U���+e�z�&�=�*�8�PJ��=#EA7Ja�E�~Z�F�0	��x�����7�,�)���N�� n�<��w!���s���W��uuum�+��JΙ&sn��,b�n}I57�_�w4T[�.���C�,|���_�D�+wz�*��Ȝ��R�4:����W�X�� �/�oP����,�i3j��U�;�Uړ	/�=�+W�Jڱs?N�5Ɩ�Z�W�!��I���mD�Y%��,��f�PGL=%�P�oO$(x���m��ᑜ*���9��:��	su��)m�ſ\��i��L��5���� �,�@ �jO�xiq�+�5�;Ɛ�^�(u� ����-	�������(jh�M�C�!7�V<��I"\�r�������I}��z�v�������}d��cVA���|�(��^jb|��H���T�%D�VqeQt·4�|N_2--�N�d�-�'�$y�pF�ʞ��q�nEI)44�@�3�}�4��6|��ڟ�(�T��D橻�m,�4t�w\W��@�!(���b�\Bݣ�t�6��#�Ԕ�W�a��+�0�wa���\�1~Ok^-�}i������ݡ�O)����bE3�>����=��Tʷ�������l���#�[Щ���r�x���{���"*��+dF�}#b@�Q�'���9)GUBLtb���Γw��c�8�JP�$F%�|���PҞ^'4�;̓F�������~\��T���
����R:�?�ڤ���%>#O2,�殍�v���+O��5?�υyh	/��w�_�[�⡛����Ax���(j�@��lP�[X�;=Ĕ.J�n��P!��v9X�u��W���1dh:Ἔ�g�3�[a�u�	`]��_���4)L��3���l#��/��A�m.ɂٸ�P�ɋ��h$�m|�i�v� �Α_�8���0ZQØz��N�9��1������?�1�TX����g�B<ǌ9�Pͤy%�d:`d���C��g4F֖�]3��/;��|n4��z�׽Y~N�]�/�(9��N9a��ԪƁd\���'����kV���J��z���/�$߶�4��"�m��@w�Kt�C�5����Mt$�=�	�Q�edd,_�������6��Ww��T��y�4�� �%޺�k��ш�m�f3q�b5����0��� KЖ�ہ��=С2��GI�,�l���A�w�igl�����}�#�s�D��N��"�M��.�`=��7��x�
|'��S�^	��VF�(���L-�*��}���r$��dJ%�vz=�����b�LZR5�p.�
���E���$�}�����-��O�a�Y���i�,���gf/{.�{2��<J���������R��Q
m�o6����+rؠ���(R�a-����������|�D��nD!��4��j�|!�\y����$P4�ps�p7Z��)�weee؛Pȅ��N�>f�h��M)�vp��Xi>{?���K�^�X����>�]����'�*�o�n�\�AE���K�9�R9f��~�pbG��gj�ccc�}222;�S��R��7h�pv�W�l�`�z ��=�B��(a�:��u�����͵7	�Sk
37��&�!��0��H��۷�Y�t1J{�W!�����ڨ�D�LU_{;	�z.dv.7�ibB�hZ�͛7!����LE�:���E�J���4�[J��w�����5�pvw���4ɐ~�4�b�k���N0�jJHK�e�j�0O}���e��4t�-)���(�d�m���![���s�e��P�uj�Nk��f��A�\{fwO�����T��Ƙ� ?6�c��G<,?	�2���CA��>����]�QMG����"^��
笠n'��������s�v�kz�j�fbb�s��H}$6�h���]�w^|e*ԙF_&�x�W�?�m~R�x�e���!���)������Wmb�F+���b��a3R��=������썞���L�d�$a��M�5�H�pq�v��LvjB$���Z��+��vTVU�>ݝ��>*�f�F����G�),zZ�ѷy.����AkX)�������|�~1�]���ߜE�#�w�,El�i ��<UX�zr:c��M��=i��2�7��!�顫��6m�������3�vF�m��U��5�
������w�X�>�,��&9��t�z�Ӵ3rg����vBfM0!-��i���&����J;�ƆJ�ƅ��;`VЋ���?	ݙ��6��}G�s�F܏�U\94��Z?K}a:#W+��Pu��b�٧����F���A�	s;����XI"�J�,`+�q�PT�d#42��³�&ub¯�?O)]�a�{�Z.�C��T�{��pl�����4� ��z��/M
���~��
���|�ֻ��� �l�)��]�._�Ltwu�NTr�tr���?+a��o��KVR��bҼ�?�z)eO6���V��Z����൫���� ��&i�If��.��C����f\Ϊv�	-��,X��J��XrD��6_@�:�M4�D�/\J2=�����K�u��s����X�6
�����������@=݄�B+0P:�z�R5�pu��c)�s����ˉ��G�m��~f�Ni�v��#S��T�$�zL�6�� �U�7�dfMMM㚫����T�9��Wz�x2�)��]�����V@��%֢K� �ǀB�
���՝�K�ma�b%�}
&��s�0M朡n��| ��>}�777��V�Aq���&��Ǐ~�Y]�n�6�.����BQM��Ho�N��}	]l�@Y�]]��xY��5`N*�-�����e#�� u��A���`K����4v�K���F��*�����D��˂��g}���x��m��@ꈻ���E:�"�'a��S����$�y�8n���Bk�u��1�դg�?̫��%U�}r*��X�ø��Bu��F1!0*���3~c8c��A��=��>::����/qu��X��y:ő��O���? 09.�����<t�����gyB��G��>u����N��,�*�N���KT�g�3T-�g��������W��L&���=4D�}�.����S���0*�A�O����|Y�W��f�Y�C/s��AVEV]Q޺���-̜>)�J{�#��_'�:�uv�nnI��;�hc�����s�'����� M_Q��6G�����2�-"��S�oa�ܽ�'�xP��[]��@��9��W{��LI���&����b��3	���wї�O���۹O��ߝ�{U�R����:�sϰ �7~m�_��n�X���i&�}Qi��R����XD?���y] �g`q$������8�(�>�u��aŬ��F��+�}R��`̍�0Ѕ6O�����իG��*_T2P�S[0�� ��m����vM��g�N�ڗ�����5K�4���r�k�t���6�z ��_�JY���i�)pM���Bۑ�nV�y��e,O�������,�n#z��Dk,�.*��io��̓�'T ��Z�F\�Α�Y��}A���?��5�g�����G���>&?�/y��{I�nC_K�C���m� ��wyys�����@oqIl%Y��'�I,H�w�9V�∪�O�^����\�}���G���t�0��)(�6`o�Em��Y�f����Nx�����4D���
�!�|��F{/*�[A`��+�#
}&��o8�?Ν��܆v;�ura����j C(�1�K�$�$�UzF�7���HF�0�(5�-�%فn4fz�mR��v����C!A��m����`��+�Ϟp'�Jt��
�d�ީ��?�����6
��l��Qj~�'�'�u�>�9��i7��O~-[X|�:b���Lz����7Bm}�J[uu�#�vB�0`��ގm."<A�����E��^��S=N�ߜ�I�fY�$�h�Vb|������j�q�|D������W�&��7��C���U�xX �m���Z�R�q���ŋs���F �o��@g������͍�>\�D|̳�r�v I���/ҷ��h�V�D&��'�B��:>!��G�|��͓�<Y������$'����5p8_�<�Rˁ*Y�lr���©N����^�wd���(�^NoQ�F�$PR"�ϡ_fwk�D>���{������K2G�D�IT/��sh���4D��H9��+/�JH�����"?��Qz��K�fD�1�u��2�����ӸCLN?��{��l�-\� �UʧqvϞ���# �觷���{R�+��_*x{�D9���DnyL ��Y	�\�Л���ԁI,e"�<}�D�����3�����}�=;ru|az`2.)ieapp�=���V蔿=W7��#}��r��h��&�������m����x!���d�&i��&���L��+-��A�O�-�\d�P�-):_x�J��͗�yw,ŕ111���,��d��]/�_���l�#dfe��(���/\�7w�B�=��8(*�I�5�4v-�F�%���#�w�z�ҿ���C�SP�����Ϧ�U���hsb�az��@%��H��Q��Ѷ�"�Zn*r�-��3���n�L�?-v�
��˟��5ꩃrBF����T�����Ν���ݥ�&�w�z#���^�`��2I �n{����ϧ��3�j��Ͱċ�A��K�ɿ��"wZW���!�>�vӌ��p�힁���������뎔�9Ӗ��n��?
*"�.���Ǐ�f�<�����Sq��8X#|K۔)V|47IK�����"�������ù��I���ߊ���<��5b����}��]O�^��QefɊ�ܦ7��,��=b�.�X}�������ɅYi�٫^�r#��H���	�8�jS�!��+!��`m�ddP�mQ��v���{���%'#��ΌI�b�qJy�����׆�}�D?G��n�hf.qu+�W�3���O�<㪢���aޗI ��ɛAk��Uk�a�n��F�x�r��M����? ��,��Lꫣ �b�}rOL��5Ð�aX\oO�G߂N��"��>Y�/�P ��=޴��CZ���xkp1�D,8U=�FR_��������
k�ۯy���¶ˢ�m,^��R������b�>���cy>�얤�=�\Ǯ�r^u���!�I��<]㟐��A�^���;\B�1���rz_SS�ι�%mܾ�	t{[P���gL.�M9��{_dK9g?K��VZ�`w��T�'�,��Va3�' `���龳�Ȉ������y������2rAW��氉H�ݗ6�L�y�>�|�KDF\삤9�nZά��r�roc3� ⋳�aaa7�a�M���"���ߘ9��,��"�;�)����%-O�hmm-IK�@�~VD���$��R8��d�d���3���勝o���"������dB
 �2w�n�6�]�*��@i���_�~9�>}^B��$on�i� Ž�xqVr��+���s����a����!����W���1V/�R��P��)o��s�\IC:��΄\��9�<@���:)4㱕Q�]��i}}R��.wff��"�,8ωv\>4������,�E�i�R�_�,���f~�a@2@�!jsW�VM��C��b	Zr�ut�A���FJ���C�<��B��
�.����ǫi7�۾y9 o��� Tzc��H���Оu*�_������$f�ȩK� ���?@7��>98�Y�6"|�4���
��zn���2�}��YȰ� �f.d�Οkՠ��vy+�>�+�]l#o�F	�
axh��C�Vs�q<��S�F́�.���杌qF+:v�A�jb��4�A����-Dٴ�i$ͧ�P[�D���������g�ك�7�}���J�W��D���jލ���-vsy!9���B��mSoN�!��|�,�~l��ɋ�XEH���ȇ�牙��Q�ǋpmZr0'''����&�+U2��99����O*����m��� K�۝�o7�x;r �����6��ɽB�/8����C���-\J��S&h��(�4uww����(A�y���t�ģ	����)����u���(�"�5�����2�0�zrкw��ŒL�_(C��x�FB�PK�ܹ�Z�����5Q<���T!!!&ox���T��ȃ���s�{�Gq��l,
S���M(�m���%j�ح���Z�oC�Ȣ��'+[�q��L$T�|D� �§�f?��+�)�S�y��Oz���P��rA��g0k����#����g�t���;@�	r��p����ae�I�*��r���
F[*��\G��Oޑ�(2��~ �~?nY��X�AQՓ�����ŴJ�Ae3��\Csss?xhߐ�2Kz�Ei���H��翧������m� �7�X�n�Þ��YK ?*���#�/��.���$*1��Dn�a�	���!�Y�2Ɨ�hJ���(EZ��夰9ҹd0@���c8� �=�Ʉ_�������L ���<99� � �1�m���S3o [�ڈ��y
)w�i4�;A�����y���E���7hIjc4�����B�����u�>��4��a�7�0�Rے_ul2��
����Ͻr��O0�tv~C]��iL�9�p��d��=� |ҎCn�z����ʯ�Ku{	����3ݗ� ݟ/�XU�B�'���n��� U�p��*�]A{�@ݦ��Β�1ǏW��7,`vl1��m�a���S��������f�<�9]}}"H�KLӟ��%�AD<@��҂�e�S����/��w2�?�>q�l�hmm�U?xpV�`�lA�-�
�>��A�}[��ks��-�%�f^�"[����}|����,�d��db��5���Q�"���9�qh�h>'�����7�l��0�yW�M�8=�ʀ����%��q�prDW�%�c�"GV��n�az^�S>c$$$�c-�V4�??E�����ʊ
����J���c �����!}�⹕O�e��=��J�������P�����Ǚe=��_�~��®M�L��~�������`�}�g�!�2G��5�����{�w@�y9:RLѓ�g1�xaD̛@���M�KHH������4������;�|��ۡ|�vd�y�d\h������.�Ԫk��R<� ��A���([�+�f��0餴����w�n0}���K}��<)����)��ME�����{u~%�0�ߴߡ'�=!��e��U���N@o�A��ӷ�Y��
@z �5�M�� Pe|C7��I���D��YB�gqi��{����?K���_ ��C����?��a���0��`�sD�6���I<��F�d�"�ws�����G��>�X����0:���1�芆��6�j��;"��sc��pG�W]��:I��$����<߼LB�m6S` R 
�yϦu����N~]+��J�C4�bv�]�ߎ
��`4x_���%J�4��r��=�����z�Vj�J��"��ʕ��j7 ��=�!��R�}�'����U��y�pqӨ����4���w�0������+�� 1(en(ʙ[�� L�N����z�u1D���w2��n{��*��C�.��a� #����NrH�i,��>�`�2�P���|5�z����K��ECt%�"���9^а�Q̡�������� �"C�����`5�0�9��I��X=$H�yD뚑h�K�M����X���0@%luu����5��C�$��N��=�ʛYWEs��.<�� f3 r�h%�:"��0d�yu~���̪�_@sh��_*�B�������I�!�ܞ�ۃ�<�V����.�C�#ȗ/]Z���}���蝍�"œ3��I��!�쉾ïE�����m�0�P@1��g���<rd�=��c�p���{��+4��K�ݶ*m�'it� 7P�$z�!����L��x����Ƚ�_ׇD���Wٰ*� aZ�O�VeC��˪&0���Z!9��[J�i]]�\`V`V��iG�z�U�ly'S��>�G��I�(��L~Q�^BQ��K.�r�:���B�����M."k�XzK�'-}�b<5t�{��vUt��d~r[�V#mo�_uQV�AJ�bs� �n� ����9HEY�����m�>7��I��.�X��~r��b�������C�9q=g�Tx�n�[�������W瘚!�$Bڜ=���o�B�R�`!� t��s!��Ͻ �΀��2�'�h	�F�Ɓ�MK�âEi��>ri�i�i��3�J.�y��t,M---E2��8�/ �'����xe�Q�z~�.<�
3J��b��P�4l7��jʊ���_��g�o�v��\}kNT\
�JeT{�rM���/m*�TY�o��s� ��@C�P����bt�5��|LXE�
s�e��o90�&��!�H�.�/�\Ho!Ĝ���J��d�rP�467g�;%W���&�Z�X�b�2߼�{g�^�N8��激��[~�NLL6�;�~��Om�'��0�}�^X1˾�p{CQ�Un����m�D����/��?����}}=������6E�Z�@���*@����8�u����TQE!SȈ�O��Ulz*��͍Oo�ܽi]?>@]��]3RD_��pォ)�=V�����pߗ���)W��gmh�Ԩ]u�1wU{�.��T�J�"�P��N�"�Ko)#��(�.~l`��� � %(F$��j�(���h��ס���������9����d�O*�8�D��O��Q	�c�{�����lyPܨ�oU��[�^�Ԭ,27��,��<�w��.Y�dRhb��(u��"6ɻ�%�\��@���K3 �Z��R��SN��q�+�{$'�.k�
�\^�{y����	���:޷�	H�e�rL;��D��3z���N�����x�6�< ß>�6,n�p�ܞ���3288H�%���;Y���I1��r9d�Cz��}�:p~�\Ԓ�5,��
�Ld�	�0%�R��a���9����R_PN{��_0F��U�U�	�jܗ�&|��z�pܳ8��P/u��_��� <Odj�����'%$�5� ���kU�șq{�&���ͱ)��7\�}�p��I� �h���k���P���? �0�U�����}�re�Fa�[�����Ew��Ukp��y�:��0ԯ=3����	�*c;PY@��&d/b�P�/�*/Z@{�?m�Gϟi�;p^ ����0�7����_���-r�k>��Y�u�Kj�Փ��+@�~����C��WZZV�1٘)���G���谂�b<FCbՋ�fEI���C�:�� JM��	�'���w��ע	oG7�K8 &R��*-Q/������1��A�dNI��A`n�o�I����"�.�G��Q���b&�l�=NM?��������>7�:�Z�����l���.rB�[��Cb�P#���#�؎�w�$Ԑ]�J&y��B�ʔo[�u���2�_�+	�W�����~�CcH"��}
/[F�����3ZW̲hT���c��!	L������Χ�8����R�����t�ӎ;v��1�RD?� �r�Sl�����8��x�9�����tP�M�>B���� ����I̒��5���8�[F��`Β�S ;�ZUy�������r�D�ߩ����:)�NxE]�8�ɃB��ݟD����-�����<f��
�ʚ
�#��&�e�8��#�?=q����&���4H�'m4�)Ed�O�gNG	�>%��ٿ@D����Iּ����Q��d<����v�c���E�c���i���ifY?f�C���9XE6�o�R2�Ѩn�M;��s����Y��� )0���=#��9�ʓ�pcS�h-<HgY_o�FU/�A�4�u��i ��w�O�@�5Q<I�vy��0C�2�H���<�g�XL���ܚ<��p��$��m��t�d��u�6��3(&�]�̑	w����Y����b&_��Peؗ�=�Jo��)--�y�����H�Ul�vh�3;��:`��N�|�g�r*g��T��
Ӿ���L* �8'J�O�8[�B�E��
0�� ���N�P!m����
���W"?��D�0�H5)2���@��f�q��О|�nG�D��������$>ޗa��C�\�b�ъ)��0����~�_dmd���D{��cR��^=�D����#�&�����p�[��Ź�� ?�B�`П�����lϣ����]h3@p# ,�sss�����jS��*p
��v�H�ʂ�S�{J������$�Bg�	��1'g�I�3Ψ�%�78�˖�����f."���A8Zan~�z��z��z��Ja0��m�X��џ��^#���}�%�3�Dw���6	���+��m�=Q�q!�(#�S1�}����>>��d��7��l.}>�諸�њ�&�d6V_!�;�P(Scِ��mݐT�4S3�������t��d�B�܈�#�c~�f瀀 "����@���>3���/-*�z���w�_��۳�c:��mr ��)!�lV�����W���F_%$Y��D-��/���t�gE(������{�7�j���ї��������x����)&�U�����1L?|���Q�Q#�2}��ɞ�UvcO��	���{���Ԃ�{Ԣ�����(]���O9Z��=�ɻ ���W�?�ȉ������6�v�ax>i��Z)xQ���0�,없u��G���|J#�:ט�c:�|�ͦ"Uc���ۨ��}���ڙaSy;m�K"3��|@�0/S�.Ϯ��Y������<�V�뗻�f��	L�0�M������L'OG���I\�B!�VFB��a��@ʛ�f㯎�'�߿_�6��x�x�5�&/OX_ut�?�yXSW�6�>�ѶZ1N`E�`�8�d��`�BFdF� �<���jD�(ATh�Id�bEP�� �2
bd����ɉ�~���w��{�?��pv�^ý���>�lQ�i��$��~�a�H�H�r�j�N��$�9,$�D���ɾř����w׬F+o��G�����[3���4{��{�:v`s�Q$z�������f��#m3��I���Źs(J��KJvμ5��;:�����{�!�
�=�I����M�՚���x��Q����m��h��hkp���a���n �peP?�Z���sYYY�.m;?��T��q��b�����;7�����ώ���vF[�8�����:��$���U�
r�9dM����EF�������{�J��/�r�}s:&6��ь��qX�3r��uK_�h�������5=9Z>L8��Ȭ�cT�Dw2����h��������ӗ�]��ëK������;�����6�L}���mY���v������S�no���ǟ�M2L�An�&
���D��dXv�Pk��б��.-��uK�;���ۓ��[6�Q�qͿ��59��a�"xpNN~zT8	~�)�i��U��>CCL'!��G']'���>F�H������/b��}�	��e�͞�7n,M�i�!���j�	(���:��>X.Y<3��a�Q$��R衼������5:�h�ɥ�w�����9��]{�z"���CC��?�ŋ�#e���n��_� �I��X''��߲*ͷ��M�4�����������zFڡbt��-��ԸH���vf�?r��DRg�_O�k�g�#K��	�5Z��_�6�VuY��]n��w�{]��Gl�EEER)���xzg����5q<`�U�SN��4�dt�;����ӟ��6]+7�
��w�\[� �<�xxF��ٻu�ɓ'��#I��L	щ���!~ꭂ�\;/95T�����O~���37�X�"��4吴�����������"���m�K�������OY�����{/�Ժ�^g?*v��p�xy{��Mpy��7gd#����]�hv.,k(�gӹ��Ш�wlP�������'b�R�A���z,�-mw�1�A�{tt��q��=vd��JIh����X^����Hc��c&�T>�5��tS�鳛�|�'�Z� �����\�G�%4لϤ�!���@�{�����8��;�Ҭ�bC�R�$�����-���m�Z(Zy�<^�% 83~�AG���˹�Qf���_|?��l5^a�� }�oJ,��M�$r �7Z}�;9m9��7]�mX6R���9�b&s�a�o�%PQh5y�[�g�H�UG�&�%�C�k|@Q�P��}�j�������};/o��\���^��rG�g��z���(�9"#�V���Z�Mo�y��<���J�m��I��+��2h�h.��f'<�O�>o/�\J�m�D�I�?W�?Z�R��ۺ��U�!�A�./�K{%B�9��æ��(��BÊ� ��_��c&��v>�-��S�jQ�~z��uѕg�`��7`�������Ѳ%�D�� ]�t5�<��L �Ti�2̵ٍ32[��<�#������$�oqm�'�ϫ�Ҫ�P��bmH͕k8�R�S������]�頻��hY�h���ݔ�h�4��"E��q���Z���4/M��`ck� �ޅ���+w��-���L�9���Pv����?��"��뫆jk�e�k�~�GHww��//6D�%Llv*��ah���T	R��� �2%�������!���Y��[e.��^��|
nG9ѿ�H�_�B��N�-B����JhKS���gF�"�ۗH���ۺ5��z�����(�N=����l�x���䌄,hBY��c�":����j���ڮR�d��u�Qc�?�Єb����c?i]���ѹ�����s�g\���Pդ���9 8WS�9��'T���EE)x�?M��z(w�8�edݒ�HT_��4�A��b�n�����,�Ԗ�R���2 ?�+6$X�!`�C���@Q�:���!���w�(��� ���bQE��S�Uo�����.��u�w�A�/��;�F��62ԼLLb�UI�=j>��>Jrrȝ*�F(��j떟�b�y�4Լ��uQ��1o��5J2x��=��Z���J�-Gx1����L7k��k�������D!R]*�9���T�}��C�^�z�<��5ڻC!mbr��PT+��&���\�j��W��n�dZ�v���ˢ��~�(�E�n/)��yad�*���O.i��GC�TԆ��4�Ri�66wՅZ�,���u��=��ak�6Q���@�//��x�Sߜ���*v+��l���ބ�U�W�r�y2>�����/؂ |�?R��a�O6T*�^{VZ�c@s}����j�,�e�)�SPL��������y�L���E
豐�L ޑ\��[e���l�s(uV��=�Ǯ�,]�D�_��PTO�O�����Fw�B��(�
J���Bd�&����P�B9[[ۛ���A�N' 8X�İJՕU�[G����1�r��6��� ��JPX�j�VDC���@�B�9DX�I&''"w�6K�;wN�Mk���2RT�K�p ���䴹��^ͯE��/_�loȰ41v}��A.�&��$-A��:�읃��ӊw��6M���qAY_6P�O���$l��[#���ޕ���,���}|r����uW�=�yEɶ'ߥNl�8�w��Z�w�3��4=o�_����d�o2ɾ5"�e�a��j�g'�&�wn�l~2�>d΍م#=��#,���l$�ܚ�V�Ҡ�U�� c=�N[�p�Q;;���_`�H�:�MQ|��FG;��+�����L���쌹zu1BO�Ug���m�L�:�3H��Ϡ`��_~izzzl���0�:N]R6x��W^Z�U�����2��<�����Qs�w�����Q�|P�q�{�lJJ��P�l����ڊే��;+���w�����؄�| �=��,|�4A�mv8��~��{4��~�j�R���nn?�>s&a]���7��^��D2D����_0���"����7�L��H��B�s�Zą��9P��'���:���J ej=�q���ڳ+U�8'�������㯡ms��,h>�=6#/oEee����t�t��� ��;Y�����	�)����ޘ����ϟ߮;xJ��H���ciAAAFF5ǩ9���J��g����ʃ�"s�Mq�*pt�CCCȈ�N��W�7b2��+�0����X�9E(G��Oc���X&Ky ���� 7��ۗ�0���A��P�����/P� ���5���D�yc���p櫰j��y�P�)@�]�����A)���T
%�.��447�CU^�b��_�j�-��a=��Z&��
����a�4��sؖ�=0�
i�~Nc�m�
33��:c�GP��s_�j�	1$���������ROf���L�vV\V��3��,ok���b,|�~�h0ǅ����ٖ��j�=�H#*:���w��TKZ��>CU*6"�m��2 #��WSm���jpj�k��� ��&�m����^�EO��˄�1�o�y�ˏeeeG]\�Bo��3L�x�@�����PM���:8;���U�˹�G�BQgQV�lls�ȏ"w͝�񿔶:���}}e	�����B�Ag'v��.4e�%A��V%An�/�� �'&%������B
_q=w���>t�6'On;+�=��wGf����?�t��`����|��/�����f��c���3Щ���w�?�JQ�����oٲ�����Q���~MY-g�p�
�S4;�P2`�S���������>/���%%��Q|���n�"�svV��
��
ԅ�#7 �S�Y5zcc���_<��h��!���d.;s挫��"��B�+#����XQc~��֊p��������h�u�sԽ7��}l�ԍp�546�C��
Z�E�LmEQ\��.������R&��i�� ��+W�B�K��C轍��4
��eF�g\=O�w�ȅ��)��^�q(M��CyCP67���!,��{�"˜�U�6�=�G��]�_�����@X�:4��!6`��Wv���54���'��d�fdli���>�|�9�1#'G266�j�����q�q�"����z�C�r�޾+o蜤bY{�Q��k���i����=������#(���Z&!���|��ڈ�2�J ��xj�ʕ+�����]S�TJ������.\� %-��x%i�v 0����G5gfFK���Eb�ő<0�����I
$�/G�� ^[vɒ%[���P�<S�����ii���$CD	(��e�z
>������i�p����88l<}��Qk�c)SrPWI�Z���2�2����i����K�Z�9��ޖ�u�9%ӎh�*�]x4 @ыe��IT���ǐѡÕ��уy��wzM%���99��2x�5x����"��e�%��*��+��F�x+pY�`�%A���������ֶ��ు#���{F&�	�&��I�?}�P,_�rM]vժpD�P��Q P2.�}�d�UH<�DoDDԍz	�Y�cЮ�x{�v�0��-	��NP���B1���%3��I���nY4/D��[�PB�c`@	K���C��P��"N�-~H1.�+Fz&+͋Ԗ/_�ޔ玲���<�s��i���)���wRS'��ii�tx_�b�����s,c��*�j��x���[�n]���Q����ɧ#���{	�Z��`�rd"�Rh�j���u����|����!Zr����_=��s�2��			��R�ԉ����@4LfѢ�`�%�^*�X�W�J�[����yn?����om���)'��bhz�
Z�1��O�b+O�I��j�h��I�i�B*A�EC#`1��D������zFn�v�4k��g��x8�<���x����zFo�Q���uy������ݻ�'N���׷9~|`�S����Le�0�PD N��X*�A��-��1�Wo �@��E/w��M"���K���

������	���~E�|�_}AQ���!�kc1n�(vxG���d�[W�jkˢ�J�٭����<Ӕ�&�uz�nގ>f�����`���_�A@N���e��**o��P��\K�$mG@f��Z�������1m�O����ً��j�]�^�&��q[��K�-�Qύ�=��Fb���&��ޫ@���+{�����F��1әj���rI!��ޔ�1�������-}�wo�B�=iZ��Wz>?i��]u���T{p��cG(��,SD��z�� zN�`���%p�P�B����a�Yש1�x��o�*c���dZh;C����MN�l�ܹ��nZ.�Mٸw��3c� �y��}���f��+��q`2G�ׅ�$�����>����p����
�������!V�_�xQ�_Z2#��>���1��eY-}4O���YV��u��8�*�n��3��b�^6;�,��XҸ�}u�����L���$����3�OK�q������Z�	SN�Kj��͌:X!�]?���r�-�B��,�<w3fS��{+o�;&�z���P�K��d�;kr��S-�̭�{h�\�K�vKz�Wʡɒ�kb-�nh-�ܹs��ڛT���x�%�D ����k�\��bQ�Eu��ES���:f�৫�����n����#�[��M`��m3���Q��VP#��ɼ����f����8�\ӑH�����@���n��!`b���������4���ETg�R�x�<�{��F�v�?�2�h�U�۸{]���t�����/�t<��,�^3�Y�7�0^���x�k�FV)u'���}ҳE��mv� ���{@Z�t���:��4%�X����Co�@/��B�{,z3f�{���L�NF���>�&��m��]�Zp�������AE�c�����$�x�4�����<�kXE��·C̺}�^�RhnԩK�'uܕ�����l���3��?��(Ċ	�f��u5�	��)��]�:�b������
�&hU���,٘��<�Ӆ~'���b��xF�&���"�fb"�ewo�i���on��'k-[��?.Z.��1�>�:�����q`i�!;v�N}�!����k �86����~{����̺��r*����Afݎ�u���EW�\)Ki!�l|���!J�˜�q���~�;$Kzf2Ug˧��\7׈>�:��^S*����M��j�w��JX��� Y���ؘ��ð?����+�$(���v(��g�+B��z�����_.~���○_.~���○�]�l��<�p_.~�����&ǂ?�ƿ
�W��X!�|xQ�W�/��|���˧/��|���˧/��|���˧/��|���˧/��|���SHCސB�`����ݹz��&��w>^��|�-��Wت��N�Ν�=j�V��),�n)��9�t����[�Q�ϩ]_��8,����_5^��=f�M·֡?�^�ݓ�7�v^��r{���oߢ�?Gӄ�����(�{��z�T���/���R�������������I��'� � U�`ݶ�������~�杰�q3���Ʒ�j��g.�Ő���l[��қ�|��!��C]]y�=<F��7�B����B��/�吪*-��"�������$� %i��6������|��-�I��4G��-=�Iڈ�
wʙ{����.O�r:h��9>M� R,�v7Au!���?�e�#𦯵�翺yY�u����?ۺ˫@Qd�σ3tBΘ�>�����_��i{9�&�9�r�5�\^�Q;Z�h��[��:�">��*��C�^R&!+�f@}�E�9B��ϒ����I4�������?��������:�
݁�E����'Hy]Z�uNQ"HqK�O��W����"%�u�h.k>y�Mj�x���;����3;�7���M��`��{��k�T��!��- ��uujτ/!�C�XdZ�<~�vH�=kw	|��E[|��/��Z<�R����b�H�tCbӝ}��1SwA^?���g�l�ӄ�gE���t�]K���N��ލ�ݻW{�*4�_�������~�������^x5��a��b���K�#��FdL3j����N|�w�p��0���z沃������m��y�{M��~b��9�*El]�g v�	|�׊����\O~�.1��S�ߩ	��|��*M�b�M�ޞ]�0#���g1���?44$q۶���z�q�֭[�%`Q��V��
���G���bQ�
�ñg����1RNJJJZ-ŏp�K����!c�I�8%�ڮ��������Еb�|!��^'ш���>48�c����9$���v�Fm����J��w@S|��������鯲����	FEPq1�3(��7e�`M_�6���}�����}�}���>�z�����LjP��hA����2��{Q`��SRS���K7p���job%^Y*��Ou��Q;����o��W/�W�z���c���G�R��Əa�6]A
]��@���+��Ж'� �d6_b�B��8��%��8v옾���(D���]�Y�`36�M��MॶLd��+��wy=+@֖��������sZ%�.��Q���Y�����?�< kS&�!A1sI��7?����mXPI�~&�N�6���_"�'���W��%d�$b�Ow�2�ד�َV�q�*=��p48*������~s� B�["8Z[LL�X�P�����T�kE�I�XZ��K�]��v,P�i�Xd���jv�M_�M._.)��X�^�2#�4h�#.9��z�*�e�_��0��/��E��i}�T���^#�:�ho�X��o��Q|�l�+,�z�C2�WQ����h�~T�q���®��~�:���]��,�M�{/���e;��,�w>|�LصClW��`�0�"96��S_UD�� N�ӂ������Z!�j8 #d��-��8���?�ˏ?ϼ2w�+Ne�֡��TH��h�`�Ka�cc�5�� ^�6y���嫒�nv�B���<wx��Ŭ��\�������-v�;�z���d�.YH6璂a�&�E$�+��w����rW�q�L��ܷ����h�u��2,,��F�Ɠ�s"���k���֑f�M�Y�#1�~�Yݿ�aI�y��n��z����Qm���7�8��p�ޝ
���!z�$�˖&t8!ҡ�v�BJȷَ�g	�m�F{X�
�������m$���ߞw��7~JJ�$�����V2�uw8C��lֻ8&��b���"��CNt���.fu��YU[{�<��������s{웝F��x�ʑAud:�]�(�:�����s9�S�A��%�1x+��ա�x���'�O��u���Ѻ�+:��.\�c�Ĉ�����K�E�:���"���M�w8	�K����L����#�1BH^FC�`��fvcoK.��3B�ޣ"�$���C��������I�C��t���zp�������zSzvI������!GHQ��*����ڔͰlV��%r��*Q����j̠�#�L�r�e*�1O�1OԢ�5�a�U{d���D�\pNd��C��H�+N��9�Yw����"u��	CJ�ur�ѫ�n��B���.{�'����l�(�V���G�p8J��L����c��dait�v]��?ڧ��� >Ml?y��l����v���-�و>�	�NK���Q3f�>b�C�r�`)м6��1=���	��;����K	o���n#}��ź�:m:m��v8;4z�kK�����%}��>��e':6/�������`�DO�B����-L�R8H��k�86D6�jұQK���<)�� ��n�e��M��^�J�������O~�z�c�Q%h܀��W�S�=C�*ۻ��߈>�	�:�&Կ�Ʀ����w�L����V(�L���̞w'bR�%����]0�ӧO7E[x�J�i�.��}ߜ��[��!�߂c���D�s�%���7u��i����(i�ouy��x�X.(����ˣ5�/;�J&���ry���l�qn"��`���5�'�㝰#��Jƻu~s���{_��z�Y�e�LD9Si����Lv�
���W�%��aH֐$�_\}NCz���߰&������հF���N�@��YE��ty$�ꋲK��
�_Z�����nXD�8���M�t S�}��F/5���i<t���*��Y�?L&�6:F)�|�� ؼ��(�� .�t�K 9剚���Oq&��#��"i0�cD�B	,�%*�~s(^6�����6A�)��m��s�<��	Y�����:���)����q�����v �x:m$��$����6�1��<�A'�_�|��ZK~��i�v��R�\UB4�kI������ۍ	��{Ж��9���gn�sA]��-Mٽ�7	����No^�-0�qƏI�KZ�F��
�ۇ�ޢ��Ĳ۳/O��;�&͝i}��S��3駺k��/�*(�<4���P�Zɹy3L��+���0�޺mυ��9����|��,Nյ��3���i�0����4�Y����w�%M�u�1*R�0�0��Ǣ�޽{���!�$Ϝ��@-��nt��I��؊�FJB<¿�h4�ƭC�5N�k.H������	�������b%��ܸrc&�&�q24��� �
s!9fC�s��*��j;4��i��@�����ʊ\���9*�Y
qt��F��%	CJ���N-]���,YB�S��r&��5���ڗ/_jeܿ?����}2���i��I0��������$���4B�yA[��w��p���':ke�\�޼~�>��.��MB��� ű��w3��R+"j�/�{31���{@ӓ��
\3y%��	}�w��j��h'W��+��PN>z�H�`�-"~���?q�]�����w�z��j�"�d��znTpc�8Z��;��L��+�$;cL��ǯAk���H,I6lG�i�C"&�PW�����]	ۯAF��_wx'�q� ���d��j�B�)�eA�h�tZ�d38��Qq#۱�n���4�i���N2�]�Z�}��'�y<A��C8�0=�.�嫞�Ç���Kn�p��F�Q�6?A������Jr����v�~���@��l%n�TE��Ũ�G$�=(�v�CMM�/� |k�E�}|wӻz�L�gR�S�EV${��1�Nл��r~��K�����_ze��ݗi�,dƍ��l�k�	�ȝ����)��i�?@h��4Ӹ��'y�v��MM��ٙ��S�d	h����c���i]���j�ˉ�������A^NɢԘmD���(���D��EZ����>�����X��8�*�ᑀ��ޕ�[i��\v,���`~�~���.����/Bͅ�cmE�QK��Zl��`r�[��5��g?61*��Ba�Yl� 2��<6�ei_g����V˸~d��H���}drz�;�e���G;��&!�<R�{P�y��<��.ȼ��p���N��{Z�d��R�D�(��z�ѻ�f;��poL��G�+���Aiw��Uvo D�R��2&��!L�S[ѓ��p���J*��ǜyZ����urZ]�n!Z̏�d~!�}3�ۊ6���P�-nVb�H��^�`P���FR������ׯW���!�$"��Y+Jۮ��z�����Bi?�=�3}hk٨c��UG;�1�7�2����C��i,�K�» !��!Ӹ�l��&�V�&���T�"����nU�֊rɾ8'�/���9�p�I�yML�삤�tٍ����X\��]y���C� .//��[8���3�Z �4F�DY�29�˨@��R���~�/�v��B$r�Fj％�c{�]{�5���!��0�ג��Mh�&�D���3SLk� ���F�7�3��P�W������8y;O�������n''m62��Ԟh��=�)�Iu�cED���꯳�
��c	��IS������,�U����f|�v�l�;�XG'r>���F�VT-��Y�Cm�J+`����x�G���Zx��x�Q�AsFz�@���H�}��˞,�Xkd6��D���y�E���*�ԑ�'j���J����&��hn�BJX�.�	0RO��M*���uE�i��P�g�:le=r�u�#�ni'g(�1;ژ�Y�~f	bE×�V455=a����N:�Xi���Y�=��pʐPft0333s,���v")�v��iUU�>�r��.[=~amz��tAἁ��Fe��3
Q�F����Y}�t��3�qsP|���k߲֝����c9��}�iWd�qW܋��>ZDV�g�쪯e�k~B;�+�c���d^V	����G;�ʙY��		_��W���Y`d��M��T��T�����*KX�Q��w�3=m�;���.�޼iS�$��Q��mȝg����p�B���r�8��t�A�I�.[(�1��.�GFp�1�3F�o�o��y�����WL[_<V��ڳ�CJu'ù�8-��"�I���p**&�PP�[@Z݈�d�� ��o�?N�z����{�ky�w\����'jV���L.�xد�=�32S�/d���!�#�]�챀�~�ظߡ��"��!#$���%��g�<������hoIl���������+�&�;tZ`aj�&�*}9��N�N��	Z����	Ov�1�I��7^�k�
�Wډ�h�z�wb���n'�˝��^�tZ\�-�^_%����+��r�$����%�����(����v��/�Z��!X����	�r�Q'�*����ۈ,K��_b���d�]����F����lR?R����1e��7]Y��:4�ot��co%|s����<
C��$��܂ſm��������|������B�8����,徖:�煝����������ӃA�p������D�S|�;�D|eψdapSk��I�ȝ:���:M���c��]qP�����	A(�⸲i�@(��s��L�;���ߦ#2D�zڻD'��M��ˮ�y`��{c�Wճ��z�
���(2%S��Jl{g�kE��O��E�+:<��aKC��U��0�l0y�`��y��p�Dfuͽ���s$O�Z��)}�Ԟ:择�\���i�KǇo��0�hTDB}ϴ��9V�������IE��AD�!K�g�j�@�£�r��$�!����cI�|�#NP.�����~��,^)W���̠%r[�[ᔾyx&x�\�Fx-Ӌ�g"�B�ĊZg��v��/<5O��RT����
g��)؋���N��V��0m3L�?����9��:�k����J��~�t��r3w!@w~%�e��x�]1*H<��bv��9��~�o�����q�1N�] �2ΐ�^p�ҟ%����Uuj(�B�DCI:���wF�=��}ѽ�V�*�;_+������?~��-�D~_��_r��޶�♈ C����ُ�5k/��&#�����C��a3vװ(���އ�^�Ȳ���D����)$�y�N=�c��"��cG\k8k�X�\�&�B��K��Ђg�-��c���r��~�K��J<S�g���:Q��Rsz9C�W��SO�#�N-&`y����OD��X��U����e��C��.�)ii��u��Q�^`��<����a��dB���뙰r(�e�C��h.++C�ύ$��4K�u�L�]��vE�!�4gtr:M��]<�mC���bj�%R�s�����8Y�Z����!6����O��q.6޳<�gb:��l�V�2�Lf?�U�<+�����V�q��w碚Nʐ�6j�Xc�x�� -����;LLG�D�{U89�&g�����c�N4�VTT<$"�Rd땐˼uK{��i�s�����a,�yJ��N(��Qv��2-Ea���j�i"�2r{��T�r�RĢRf��z*�:�1�y�!2d֡)@����U�ȼ;M����\�/�
��R�F��0w�[��U<ގ��33�������*�.��bټ�5?��x}��d�!~��=����ZȐUnР�J@����CD�+6G���n�͗N9V��ޗ�1�$�Y�`�U�8�x����gW�Yb����B��QI��.��F ^7i,3�}�t�!��<-с�}[��J��S��#VM��K��2��a�ݑ#o�ހ
�'�����8��]s�ξ�76�gg���N�|��S��K�O ��o�=W�\魼H�U@���y��~y`���F]�L:l%�2V{�$K}��u���P��N�A���+-�����������i������֒�&v��tP	�@�p�M������ڣ��\v���w�<-�/G�$mO�|(u���>�ܟ��3�6�S����w7"���d��i(���/݋������kll,��ZԊ��U�S��p���T�4EU�?j�� J��ѦNv����֦��Y����WeO�i�k;����k�����(�jPI'>�v� i�gh/��w#z	��=x�,]àaH�V�]���_�������T!δ.GI��"���Lt�!�ۡ��y�9��PBKT�I�xZ�6�Ȋ�k�@���`�`���N��%�cl�����C�VrE�����Q�&9��ۼ�	v�Il���{%��q�nk%G�u�ʪu	����#Tc�\K]�h4&��_I~��/�W�ASAN��v('�����oe��~�
1뢭��e��A�H0�=�z���l.\^�� �t�%����@��� ���[2O֧��y�f���t=9�Ξ��h�RgD�1�i\�p��XȌB6�S�.)��x�tK������GԄ�sO=�/6�-��}�+K�"�ڇ��?p��k���̍ı�����?�̑2��~찑�\OUi����d|����c�S��U5�u�]0Wq��|r�,�7�~b�Lò�E�❮��港G4�TE�n���,���/4��~�Z��sӴ=�?S��V|�i�Y �?8C-($k7r��FFFVJH�\!��� �P"�Ÿ^���ר1�I��j��A'��Y�Q ����Ij��?C3���)m�F|�&q���sO%E�間���W�2���b�s��%5�UCS���1�*����}5�&����D�+�Fw(?�^"=���gտ��4F��5���ҽ�N�9��I��m�|II��2%�O�ٍ�;�޽-�Qi��Oΐ���OU��u�p����=����o�!ghH^kL�r��R�%IXp��<�����!�O�+�X�i��Z70`n��Y�66�&Z�	.B�Y�3����*h��0F������ϱ�7�|�[��6�n�4v�y��b�t����Dʡuy�2l�l�K�a�܇����`��>�G�z��k��3 *��-����wN�($�|L�y0�v|�]S����K��X|dH�a~s�j��kbX�Ӫ����C1abĸ�"�o9��_���V`W�:J,I�>�M�$���ơ,m���Lï4N$���z?L��\�X�gv������� �I�SG��H�|���(�쀪ТV9���X'�Ơ�����5挲��Au�Zr�ZR���yv�Y���[�T\v%�	��&�>�e"��ZQ����XY�(������fS��*n�.�"�Eh^*����(=MWptphҒ^���Z�y�7��^���X��CY�X��0��F�C�dp�j�@
��1�=�%�ɒ����gN9���W�c�cIL洛��	rJ���f���U��4��8|�gA�q";uR��M�}���M���{OU.��%�C����uu�q��=%��t�w	��*ӮZxf�|�V;w)5Mj�\m��s�q�d�~i��7�3��[ڊ�~u�����&�v U�E k��9b�@�}��h�����=*g�'e�=�6�4��@�����2�944�oab��Ig���I��i��z�2�b���L�SNkν{�c0����.e@s�5��$(rr�zL��h_LD���z�%�f(M�Eӝw/�c5	���ށ��ÁTW;P�;j,?��VM"o=ȭ��ق:�s�qTbELH���7y�32S��l�3eC��#J���TG�o��CC\����f��#X���m� ��%%��S{Ʊ��Ȧ�Ä�Ɇ$�����W������t�~�z��xW��%J���(�r�8��*h������ͽ�Dy�nN�t?u�q�T�&�Nk�"�P�����!�1377W��a��������}v]]]9f��H�0��G��VV��:M`����u����#4�8���)��3ќ!o�RY��m2��iP#�ac����N�u;��Y%��krVR�����9Tr��;�n�\#�vYd	�X�&�����d��-�H��p(�!�6	|�k��M�4��-���``���D�(۽�"A(�wi����ɳ��<�J=�����	���Y'S�lo��*������;��-]���Yo���Z2��M�+��Kk{FR�ъx�V�H�JN�ݻ��⭜����)�gD�|�@����"����Q�?�+��뷹\n��~����*�`d�`<����&�kG�\P��
�`#"<��yB���sqm�OE4����2�����2TY�r�Ni�B�w��o�J�?�5OFI<��s�˷�O��.���O�eT��"X�ho"��D�:��"�"f�e���L?�\�����䴨��'!qįh�|�?D[������yvc7Q��O)e��)�%�Kշ���g^�q�)A��%�$(3M���-����y�U/�yZZJJs	��XBcf���T$1Je�{d��ܘ���~6j�#(��]����������qq�°jBdI�6!�k�����qI��X�|�$�j����x���555�׎����R���=ȰV�Iy���N�_t���f�s�\���ڟ��l�7<��貖��Vԏ�	ԣw���c�6�F!W$�m����p��]�&�Wj�C���J�tel��DKօd@-q�����C���"����C���$l�b��r��[���L#X%��r9��U`�}�D����`t���(&��[ԥX2�z�CdA���	��W���)��{3�v[ٝoτ�ƃ���3D�ǜ��[����8"d��Qo_�ײ�ں���~�e_���p��8�p|����z=��[��o��}$f�pU�����Qm\��E�6`�ȠK��:�b�u�P�\��K�1G�\GnFĜ���_M(<}A*ݱ
����U��?������&օ.�By�Du����F���:o���֯�����cx�8�O� �[��P�l��C�z'�^�=QJF�D�넢 ��/���0�1�r*�S��S�����>�и������DF�-V�:F}eY�Xx�{�A���-�6:���j�j�p=��Cw�����(�5�<g�&��~�w��V��#ԟ,��n���$�K�Qȥ���{��z '%�+��zZh�d���m��h��n�Ih`��\mHp�#� ��5�O���K��ވ���,��{����r��E��	���
�!A]�H���FZ�<�o�Y�ΘQ[����y�|.��R_���t4!�Y��y��b}���ȑ7#�V��k.��[�"��r��#��%��)�kG���#bioo���^�.�:OM�7�J��DQ@�!�-j�s��%An�(1RjB��7�����$�mK�����eH�͡��lv��O��j�vF)_6˧���>TF��o�y�5�~����ˠN�;;v,���9"����[N������J�t��Ut�v��`|����N�.	�yė�B	i�'�R����̴��t���D�zW>�~�x�P(lՔZ���%!�]RF S��g�щ�ΐ�<	������H�����'��G1;]�!T���')(v��יh�*�tQ���&_��X�O{����過Y�֕2�?�;��r�djC7P5�5�(ʵ��q��?85O� �-Y��M���)�^���xH13�Ǖ�=��������؆�4nS��b8+g�o9�9�)fh#���%�[���_<��gЍ	)@�9g���)Ą� �õ��YE�갅_��Ox^ I(:
�"H�����=�ë�r퇴[��oJÏLf
�{^�^�r������<�!��Ƙ����j�JR��\1�%�~��gup7�A,b�I��K����s/V��#~�~�&p��E�#��;�i�Ԅ���#��~� �.�>��x�׽�@�y B�ie�I�����T��V��<��z9���A8�w�(6�{�ՄSOY��w%��v�=��ۼ�U�g�n��@[�?Zrܾ�"���`֩C-^+w�g�(��8�_?Frn��	�<v�tK��X:a$X=�k+&�"�����LN���Q0~Vk�/�21����5���w�ʵ+�	�7Cb�Df�Lie���'�!�Rpْ��cפ /L�5�Ί�6}��Q�u�%r���NN��萷�8¿>li9�������"�z�憦��z2��g�(kK�]�*��Y��>���H_��'�uے��#��{��S�jB��*,������c.��j��A���P�7�U��c34�_��j�Dp�u�C����@�\Ǵ���~�"THّ]�K�	G�{�����!*����)��ܽjj,�`oo�	 Zǽ��(ĨR-��»y���"�9��������i��n"�%8e�%��"%%%�qJ�o�_������P̢�~b)�9���"ەl��ty<�_i��va�[hÚ�r����~�U��������z6��y욡�˗�n�1��$� �ju� ���֒�\�.���<Ra#n�#Y#D(�I�_�N�Ԑ�N<��X�M��Rt* �ҕjVۡ�<�N���(�qC�k?K��rqee�5fG�Tr*۝��W���h ��tP�zt��x��)���32L/AA��a�[}��ک�P��@n�Q���X�8�s(y��:� ��B��goQ�đ̪d�N+�	��X����l���x�]�܏��5���@F���')>�=�����y���5�"@0�r�A� X@��i:�]�3������(��0��$�!�A�����J�3���[��~�)(&�&�6
'I�r9��<�evM��Q�����e�/_>���K����.�m��ur�U�K�S�����9�__�?\�5!�,�]�r�X�g6P���Vm�߈S�xo-��t�Vvיڍ��^�����D��jFzZ5���j8�uM
���䜈��@�1
ـQ��2��]:S�I�ѱ��ԓf��j��o"*d�\ ~r��q����j�:�s[1iH�x
>�+Q�/��ȿ��G�{(IM� �*�B6\ܻ9������V�vLN�7�������-��M�=~6�}ͳۄ�E��@����.k�*oB	�Y�,,��>�/�	�쯾3A�h� A���Dm�E'�b/g�Sܙ&=$��z�Y�,�>.j�Fn=��Ҥ\e��"�W�kį$�1��:�����)X��"tN� F��f���ꖢ ��:O��>���Z���X�r����/��^s��]��P��\�#��=�{8�i��{�$�~<�λ��7~��<d��۫O�&����e�O�G�{Q��=�u��v���U�{-��7���3��U(�9N9�v����1�"ף��	*�w��|�w�������0k�..�Y끅�!��n%��n, J"%5UKNN�ƽ4��(3'߽�ʸ����u?�u���~H�/X>���	v��N�ՒPns�'�x�;�@�AM�)�ދ 1&S��(-���,�Ă��A��k?���,��i��hg�RL�SV&�_���r��h��"v����F�y���(��i���:���rDkk`�wtoH�8����Ī���&����l�n&��~h���XD����PUy�	������ce�g��:���I��K�@�(����%�a,E̺�G-������ߠ���g��Lf���F9-Slv����yE����A��3����'�̲9Q�����Ch�_e&qZ��V�z�5��/1�����%Z�����ה�.ҍ;��>��Ri��Ҍ?ˮ1���a����>��z�@�I��T�S�+��zk�v�<yc%��3�������Q}_�mv�Rd�w�[t����5Ǩ��(��J ia�Ĭ�2�J-^�:~Q& N��i����8ik�_�֙u'�.�����5a��w��V�1�aw!{�5Hk�]1s���	�S执��?~����g4�`�L�offf�	�C�q�\�bC	�]K]n&�R\����گ�6�&IJiyw~�oyĪHCZ�M�q���:`��w�O��R<w�U�ps����V�9�������b��ݓ�ĠW�������í7.c/!$g��g�C�4���g��w�m�Lz�5W;w�;9̺D>N*$��׫u����j�X:mz,j��ɗ�a�g���Z�_v��IN�v֦\� ��_�����;��v@ʿϮ��O�d$�NNo�ѯ�B�:�s��ū�.�r�ϻGK�&�f��=(6vin{�C���f��ࣜ��M���{�7��g����������i[_�Z6(����!�5�"�E�@D�@�~�}ĉ#��3XQ@�(q4,Q�FQ��o̍>�R�7��{��{���~,���2�Ӕ����w5�j�
}��D��=�!��H��eR�R==�H�Q�/ef�?���nD����|��_Q���<��!���O����u�Ɖ"��~��:v��Α(v�U���&=��j��,\qL��)�4-qJ���`q�:z�␈��� E�
�Q	a[�l;����*\���A2�ˎ�X��N(���u6m���8��bVֈ;xZw���׏����^���θd���p7,s+�5��'%��8�U%b�8�fr33��!+�Q���[&���1���!D��K����#Ʌ�\�o��a+@[�˵�e�da�.Y	���X�ҟ�`ہ'oWh�-T���*ZNNNk��J��9����,\�Dת�(�>U�Y/r��p��4MF�=�?�|-vlԏ�U��J��!'w�J�w�Ĕc+�%��/)»8ΐ{�J  ^ 
�>F��_l;���O��:@�BZU��w��ۋ�Jm*���Օ6Μ<�t-��LƭǞɻ6�YB����X�
�c5�	>�K)�Tff��8��:��4��z���٣��@�o�lNff�K���k�\|�~���Ɓ�V4{R�MI�߸q��''����0���au�K���@�%*f��C���$��������t1�({����3����>����?�Fg#d	9��F_M2������5{y�o� o^� �ݭ{Fă�'df����V��H��Zs�\���ɠs�XK᛿x�~�w�]�C"�N]�G��-��eӣc�7�r�Y�jH�,�^�?�N�͜����!�`M��~��u����~�����Č�Bg5�3_���݇����W �����๳|w<�qi?���Gw��n&���?K�ea��ZW�L��f�k �O���+�Kܔ���sY��wtc��#�1O R�@�[G0�o��A?(��V�g���.I]t�#���[��E���L��v�&��1pk�k�z��	4��Ix�����O��V//�ALL9�
W��q�;_��U^�+M�������l������[���7�KJ�&��+|ޏ�� ���>��AV��ݹ���CD��_��v����"{ֽ�i��j�b�.z��E,��,?��
J�/���.�u�yw�\�?X��!nT�2���{�8ՃD�������D-ӐW����n��AF*�i)��lȝ�ַ�9����<<�$V:�v�JP�x�-��y���?Rec����u�_�RH�dK.Z����7�!I�H�v�����[����l[�N���]�����>���t���\�="׳�J�mҷ�޽یΠq��v�ƃ�6��c�ݤI{���Y���+�H_�u��g7��3)-���mA�J[Jcq��$Դ�k�g�����}Tԍ��Is�Q�E�^��F�e�>?בF==g9��Az2��p;�m	K�Ŗ��糥�7 �lG!���?�2��3<��`���t~����D9������l���|+��X��+�O��)`M<d��<^,�i][��	�RZ �FOP�̟|||�YWH���n�D�5JT��[!Wc��s�&v�%���gpLS__�J�]
������NG�$� �A�S�b�����u����nz�+j����Z��!�~Q(�|-�`�f�6�7�����~xH-�[Q䠦��چ]q��85[$*�I*@<d7��9#����(1����v�$0��DY��[�f6�p�b!��1��� G�M?/{�RÌ�I�Q�)���H��2���N:R���|��e�&q��n���?y�~}Bqa�Ǐn����z^~8G7B���.h��R�uFo;���f0�;"%�}H��:���E�*�����,f$F��U��7��
�u��@����%�N��O�+:21o2M;��7E�����n��n�g�u��r����v����y8��k���4������C��ʬ�&:�[�"��� y:��>� {�b"��n�]nۑ?3.$O�L�~Ȕ�O��xU^Y�c�G9��ƭ$��6���[�-�7���p��9x �U���
�������]���� "�&w�o�<$�`ڜ�����y�Ђh������
��Syi�K
&R'���Č��G+��L�m&c�-+�|�6���̧�F.=���1`���JP��¦�>I�V�av����&�����o	�U�ڎ�R��_�~��<=�@E4&C��i��p��a�j�u�y/����|>��v����iW� �𫦙�d]]4g1�k�Q�ێ���x���4���t,�~�Dq�F�t#�g���%5l�F�-��ִɊ��;T
�����Eާv^��7�x�+4r�P˔��h݅ǑCX�Dt�i$ܘ�Y�����;��j���;�<���J��1ߙ�25�7��hX�����Q�ω,�c��5��|>���G�:��{Ď�Es!�cSe�O�(�d<�]q��{䄋����.���%K�78>n7�61��qW������u���B��3 :��Ш!o�k^�ΦBfے��q�.d�3�M�M�!���ˤ!��I�L�ސ�~XM[�m2W�2�ʳ�	�O�>�F���I��b#`�
H�W����i�*�ã`��8��3].���M�9���MͰ���
��^��a���{x���.:E�;��%�P3�\l���0�I��m�1z��v��jժA�kw�r>C`p�'Y��d�|I<�������D�L��
�ƀ`0�Fz�Zm�I�+v�)����F�O`��YO�2����t5F>j�F=�P�2���(|��?Ě���6\ugG�ye�i���ш��=��"$�a6����� ��5���oY����#`�|޻p�,�oH�0J�VyG�C��sS{<x��(|�P�]:�;��b[[}6o~v%a��IW�q����O���������酹i!M�bz��L�������۰�g8m���]����
�5z�B��%��H�0����A6B���A �Y��k��r�,^=����Si��◔��q�#c1_joAmU3�'������33[V�ܾc$����)���lm�S��[�m�2g1�Qc'Ǽ��44���D���uq[R�c����Sxu�X��b�e���m@u,�m�����t�a�:�DY2�'p}��Qt.�`��J�l$5����� �;<ǅ���L�&<E�p���).���]1����FF��l��E�Y��v�4���f{���GqNGtR'·Z�`yH�-�s?r�X5�h+o*�	
���5xֺ����&���&3i��?Rv���/�����f*J�Tr$�p�E<$���au�v�t�^D�9�3�q�� �e��[�ϔ[uE~�<��(%����3&f�2�}�mSp�v��w�ܙ���9�ʁ�~E<���kܓe"���^$������^[Ϧ"g+9!�_�Z���e�12��`���z��`����6��Tf��0��A�`��P�1S����mY�z�]�$ FNsS��UHa���f�X�:���j����r4���utԫ1s`_���n5l+X|�j/q��߄���2uȣL�͚�F��0����l������q�]�a�b���&P�'~��E[�wq��	�T`��uUl���ׯ��%���R�D@�ϵ��ۖ�Ӏ�1�7&������F�m�
xS��� 8��V���y�zL$��S�0<��I�Fb�33��Uj��1Te4�(�vj�"���+3��c?�J6��W��Axq��H�Wf��Ԅ��]�.ŝ[��_�-��= ���\M%�kyE�Ak�K�������.���������&��:؝�?Lh)i�;U.�}��Y�����'�n�[�D�rO¤��6���.q��vu2.�-(��H��(��=�g�ʹ@��l���� ��L�tt�6f�'�,�~�p}5b��JJ�����tTB�[=g����Ss���Xﺉ�F�b1�`-	�uu�3���2�Z���|6b��� �=��b^�*&�N��B��<�ሒ7#˵���?�%V��ӳ<��T>l�Z|� Hј�e���kF��(em��8v5/�k͎����(y6
�3#v��D
��^͎�#j�yYYY��P�䐑R��s��
S�Ջ�U�7��[М#YmhO��gΌ�c��e� ���:�NDyY��˦MÅ�ù�\\���m��- 7mA�H�4����Yr�y���K������s
D-f��K��6	C1(5��׮�KblFn�n01�|��(%9je�6�������^%!5����X���D�+�����,ᾤ?���`>K�0�m,�s]T�K8'f��\�tZ�H���Bz�%��[�ʶA�n�c"r�< ��D�%6B��`��S��؂5��E����n�^��~�SQ�5(����ŦBC�?#��s��G�����Tnʗ�J���pu����#[�(4��Ex�]��j�D8�>³�lL�+���"�h�D����|�B�������D�X��P�������9a���n|We�F�da��+��AXm������@��_J���=1��]�[?�g��^���� �}�����.�5��=��y�n���"5ݲ/S!��}��m��kD ��}���DL�D���CeuU���kK���;����19ݥ8�@�-�˒�,�aFM�lCi�s^J��Ơ�{xk������O��<�������~4���.�DY(`s���s�Cm;1ziE{��en  v�-WZ�TZcrB�1-��`\9'��hJ������OR<�ƚ9窐����*Y�pb�E�^�z{�J�궉�u�B�9�,�_��\�}^�q�m#eo�$z�>	6PԷN�@ّ�괤��H��j�:�e�J�$X�)h�E0�8ÒF��u��Q��qZKs�xQ壝��5�WC(/OO�4F66��?{�v���N�nlf�a���1�p�4�X��ȇx����$��ppuՌ�z��H0bl�>�Q�),J���ˏ���'�Ho5Y��Bf���`[���z�mG:��D|�َRݏ0��c� �P�>�*�CL�
㊅�$]^a���t�����()��i?�iN�-��c����?~r�.E�K��� `� �$�ϟE��vA!r�2�l������j��e���^�N�M�kE��ҕ��T�YIW78�'��s]����?�-�;mؐ���E�8O[��>�b��7!�o�ݾV��յps4�cmŞ��H�ZQ5��� |!��[�;
��![�c��6PU~�8��u
�U��S��3�Wc�����x9ZZa���k��������e�����8�ۈ9�o��9��h�Y؇��uA��ӯ\�rvس�Ѹ;㳒�Z������~��ne�"f���þa/�œ�*Fg���N�e��:���;G+�����vV��ʟ~�G&8�=���z+Ȟjh�
�m`P�&ƫ��ܧZ\�{B����X�H���s��I��A2��qS�_�ό>Y�'@;S�ѝ�Gh<0�����T�8a�'ħ^�6J,�c�wx���v��n_'h���K�(�O}���aQ����;��ow@��B�D�b�q�+��P�G�޽����E��UbZ������4�z�  �^ 73�3�#�ع�7|x����F�i�`�zM3ng�eБQ�w9�CbdZ�q����~���~I��PΓ��m1��u9g�5���	��R�B�<ؑ�����H�h7��u�w~E�<�� !���$Ƌ����4���l!��jo��GSccT,{x���)O�PV�$����q��}�p�o��nᎧ�!Ğuqv����Z�����s������+�g��f��ƺ�k3w�R�� .5F�������{�"��nK��d�C���5��ëن��Twf�AᑶQ���X�Wz�Z��w�T��`*o������!�#�p`�q@��7B|����ŋ����X��6��T�Ǉ�ʅ�==�/��I�����	R]d5�~�s�S��*G�,մt��Ml,���]��Rn�i���x޻� �@��(xO�$��xC��?�
��+N>����d�F����lݹ�i,fz5�\���_���DBD�f�]����L��|)''�	�JyS	���C�B�
��|a���O&�4�a$�}��^�IQ'����J��͑�b`��GR�>�
wU����wt��p�X���4v��e5Ht��*?II��7�̶?Pz]���ll"�
h
�1oY lTg�"���95ƹ�<`�@�^;kv��^W�M\��A�3n2z�Q$�?�O�*Z�SF��7��4�֕�Sl�8���_�mt�MCv�~��{m��G4?�}�e�O��opPݤ�C�O�e顇��#�Wv��?��昋��	�_�1QD祪��?���dD�fj��t�~8����|��n��q�>���u��ٔ
L!���AGky�QY�ME�e �����砞�k}��0W{�-��XJ>�n:�<�=�p���O�QB � P��d�\��q ��F�J#[�E��P�y���%ާldz1B�.v,�_T鈎�^ɫ�������ZЋd/!�-%D�����T���;+w��&�Ֆ5�D���έ��Q���0��>�v�Þ楩$ܔ0۞�"N�֜(1E �1�ˇ}}}�A>����0T�,�!�@�v�?6��.�N��%*$�2�
���{�2�@V�;�&|�tP�h5�/k�����Բ,�D��N�z3&��������Y�������B���]$�Ի8�@8�\Z�6Q�>.��ZʴH9����Z醡�� 3z����Ӳ�aT�n��ea�..�,���=d�x�߇�_6�#��y�N�����%�5�`4�����1�j��K�=��;7�B6>^�7U����y]q�8��܆�BP��ۻC��3�!�_-@}2�$�ڥ3���&�ɖwJ5WV����7�c=��K}F�j���o�}[�D�w��7� [�r�n��/B���F���d��f���p8�����= 3�σ�o@�	d�#��Y�%�3���7\��O���u�Oָ���^mn�h���YVh/�_�
T122��ɷ��A�f��{�ғ~��m?Y�����Z��+�I,�U=K$��ϴ@c7h�B6}2�&�q;���>��w�קԓ�XZA�f�ɪ��U�ވ�#�"y%8���ぎ���l;���켼<�j��&1�`�2�oh˫��^�k\�Gf	��0h���#o��vY�u�l��3h����U�����V-`��<�_�~��e/�n7g�[�A�\��í�?�]����Y�A���i�?(q����a�d���֭�Gy�4��ڞW%�"�;D��]!�;�Ʈ؎s[E�s���婜e�Rͱe��QdJ<�����ib�f�L6��P"@����b�a���]�3'OP�� ��G�h�c�t���Q�����q&$�R��`ڌ^;�^���&ʕ�@���S<��u!��?���|5��<���5p)�?K&IT���Av�$����o�H�4%�f<�S�[��9ΚU���@����7{�K�^�Q���}��LZ���^���r$��|v�����i�j���4�s��s~��4<�[��^�7��L�>o�(CUC���9:������0\/%;��Ejj� ���0X����>>>swf�!����կxx/�3�;���P2�zHi��Z^�܌f������˗��ə�A�gO�xդ�m�~L�� gr�4�t;x\K[֠X�s�2 �:900���; 37��v�$�9���S�6�վh��+����� ���ՠ7�������2u�-�ϴ�8��a������\�ja���0�_ET��s�%Kzy���<r����R�UM�{�Ǧ�9U\�Z���D(=��q��w��/��I��!y��#�)������Wo���Uq���٢_9��?PK   ��X:�I��  �  /   images/684f3f0a-9a9f-442b-bbe3-87dc70a48100.png <@ÿ�PNG

   IHDR   ^   �   [�7@   sRGB ���    IDATx^�g�e�u&��x�=�ܜ+CYI �[���n%$aD,*PH�7zH�����m=$ �$$��L ɖe[�H� +Y�n�'����Z��F��{���FJ�N���s�5�7�9����WA��W���R���JF�o����J�+}�����g�{@�q(kH�����R�c-*�V���c5����ݴ,�R�j[�
T�Ď�$�R�I�"�mY�eY�#۱,�rl��?��X��F�\?���M,XN/��Nl;��45�I-ϲ-�J�_׀R),+�ϳ,�_�"^znj���8�)ˎ�)�4�S(����ہR;�.�ۿ���]pA��z���9������|������/� e!�@h뿇
�,��%���y/ߦl�hi��ߕ��2��_����`��=?c�=�e��Z���"�{^�r���s})�!�3\�>H�$l�[�o|��k.9�1��W��?m6Ñ���c��Q��bAԂRJ�R8r�),�bi�T4`��ϛ�m��s���+w�.�Z��Z|�~��/���GXr!�:,�p�(i�۶J-'M�ġ5�������'&���m˱-([�J�T~�Z�~�)R�XQ��p��f�_}��������o����J��\�F�o��z���MJ��I�D>�#J`;b�D�vl���m#��G����A%
��!J8��0����hle����#��9
i����Ba�u]�\Nq
��`�6���;�2�Q�m8��8��`�{|Ǖkm7�����^x[��Z���D��]G�RA��h!,�AbY�r�x�������?����{3��I�[o��؎��^��G�z��}�0�J-���h���²}�$�e!Q
/(I`N+A A�i�|;�,��s@�W���9��Jm$q+U��B�� ��T���C�E��E�V�-�D	�|ql|�J��	[�ȻlXpr�*I�~,�Je���rE�|�;W±b�.d �v�n%�<a����>l?o[�s�o~�ͷ_�ş���z���W�z.�c�
GT<�����k����	~(V���m(���sM*�s�F�ܸ�p=*I�A8�7�t8�a�%`��:HS޸m�p���t**M��n�q����x�J�������A��%Z
��vi�B�s� T�\�)\�&�`��]G�����o���O�j�ws��3X7؃+>�)5�i�>kc�C�7�^3t�?�O��&�?�w׬�����zugt��;����{P�e{h�cx��-��6h#��!��\�ڪi��j�?W�ޜ;���X.\׆�(4�(�b]�V[�=�w�r|��h�X,��j�������n�P���$
��#P.r�"f�pG�H1ڔ.�GΥEH�&���(@��<�Np],���2�T��T�1�b��n\ú�".��?��hg����#��}ޚ5��?�k��ͅG�k`�O/���]1������	����h�Xv�V�q��v�E�������y2rT" �/�ٗ_Ə{�����c��#
"x|8n�$��wN9'<�-E���v�x����ǟ���$1�q(�fs��c�yG����'�@�݆_��B#w�>�߼vH��{'W��N��N-	0�[�����F�R�\~�H�/��}��G��b�GqE����Uǆ�|�O�f��]�?����?wú?��`ͧ��9e���_ܽ���Ќ����	\��ۨ�>|��8J�}�*��BXq�{���yg��r^�&��B�������$p�<r�p�6Uǎs>�S��npK�IL�����m���w ��z"�+"g�@�B^��#��?�8�~�:4�1
EWb�����~<��s���s�
��Uܤ��6��㻶b�~nCj2ڟm ��/���;�����#�R�]���1\n���X7ZHcL<=5q���|X���g�x˹��q��uD6p�_�Uw}�$�
���}E'Eژ���N�<�4].�A��݋�>�c\��nN	�߁V���8I�5� NZ����>��� ��Cƒy8~���#������Dn�p`�Mtz	�`���3N>�(����r:y|�����@��H�$�&	r̋�El^ۇ�r�Vl�G4�Z6�B'C���*���M��9� �3�L]E�,�P��;n���X?ZN�b5������=|�?t��_qѮ�;�����o<�+��6�|7
������`�P�Y��w�s?�\҂��%�˽�ޣ�����P�=Dn��C�0gT@�B%X�,.��a|�ݧ ���r�2B���'��;���+j�l[B=.��U�PكӞ��~r7~��c�\�CD�,��T>.�~/���kh*a�Ip@w�+�ς.`˚n��Ƕc�H�FU\Mh��R|��/��N~�����"CS�j���1�������\ߟ��?>8v�kG��a[����=�;w�2七�����a\u���Js��|�:gx�����q���� �1ڵ9ٜ�J?���3�����Bۆrr0�NT
�e~#o����������A}	|��^���S����Ad���g#dk�pT���j��s�I�t쑘�8��ׁ�.�kn��z�_�B��/�j̹98q�4�i��O�>GoA�:��w��������7�Ѓ0q`������B�U1X����	l�0�����3�w�=�w����[�{��]���ϻ�����#�*�H\�a�8L$�b\5gq�{~;?���E�/Έ�����֣���ދzd�g$q �w`96� D)�>�8�=�^sJ��Εx���c?����[�0ӎ�H�n�KE�Zȩ:�����lA����Rꑃ+�|y�Y��.��-�&���c���y��O\x�uC�"{���t��<��W;$���$	:�E�v��5�M>������6D�5�����[���d5��+vﾽ;�ZzĻ��1\��{�t�������,�5q¦a���o���Gl���,^zuO�f�<�s$�����f�x9O�ٮ��q�`�s�:�y#�y�x�����L�Ǟ�5r=:���y.���g��D�?�q,6����CWw{�L.����?�+���"LSI��@��)0dѓO��q��;p����X��O<��fjx�_al���ac5�Yk�b�FԚ������Ob���dRa����{��9���O郷��{.��r+]�smg�_?����.��7Vp-	��H=;A�j���w�����Ə�z�߶Sa(�^�&7Cf���giDi��� �4��4>~�i8��S�������v�FԒ<�[D(�~`8h9�/� ��U<��;'��d�~�����/ @��C�q!�h�(�D+Zq���E��u���'��م�/�
�kP�N��>O6]�H&k�S,�H���ܟ�W>�	l\ۍ)`�῟�k�����-��o}�����b��"�����|Q�v���ka��t2�F(Z1ri��wo�������_������$��-�1�l��*�kU��<\/'7�Y	�h��\���x�o�����?Dap�[Z��B�J�l֑�y�#�n�΂�(=�s�98꘣�����C�?	'WAb���Z����y�r�S 
Z��[����	|/����1����p+~��Ax�4�r�خd�\��w+���X�Op���	��ys��c��������6�p�-�^�m�7�<{l����qãϡk�	�3aƙ�!�V1��Q�l�qk�����|U�x�)�ے�����pEc��9��i@{oݲ=]%L�����a��0ӈ�Ps,Vܐg�*�6줅��q9��7I�3=_��Ԝ$BQB"��d��+ƆcNԆ�+�dp������,`lf�R7�a(\W�m)��'Q(�ړ�!��|�|�q 3���c���;:�����7޾�3;���`�^�}�)���C|�;;��
�T�9��L�|+EҮ��E���O�_��.v<M'TXGGї��
`Yd1=�^P���a%�$;!COFvN"Z(��b� ���v$��ȓ��C�a��
�B�3�0a�-���rp��(D�L�!�h��V�� �2Z#��\�w����p�&1�����g�k�0L�tb��s��>y����-���r��)��7<�"���ܣ��l�	�����#�QB�
a�)r��<��$��<�^�1�b"�_�v��:6mI*�I/+�G[ay�E;��Z�A���	�I1�H"����rIQ$qKr�\�C�l!_,!�`!J:J%��u�V�PЊ��R�1�%��$(��nG��	�2M��EO\�a�v;�@�E��쓏���ᤑ>�(L>=9}�y����_�m�>z�_Ul�] :�<�4��/�>�xԬT/�ԂC��r�pR��H��2���9�lW���$���1�u�-Rʌ���Nʇ`Ny���41�O�֗*mݰ4�,���4yFF�[���2��,�)]�r��diI��:�-ߧ���ӽ�s��!;��I���Jc4h=�c|����0������;F���a[<���������y�kσ�b�$�?v"4��B/$�	�������o�.6^.\V�xc�X�� q�`�$��p����ۢ~������J|h
��暖^#%=��J g�N�	"?���w������7\Q����Ld�u�F�-��9�K�� N�'��~:>}������\ϸ����`�_t�X_��z�9�+��Bb;r�di��P|f�vic�.]��V)�6��E,^X:��~�ZE ,%֦A���G[���򳳲����~��,�������"+Z������>_���x5?)�X��Nc�4�:�K�z~g��>��OƧ��}d�+��x׶o������~�E�7� ��� ��>�����(�Y]9]%(GK2���� I��҇,U�W���o������=��`�Ę��\P�г�����#&,��.T@�+��؝�Xۨ#z�q\v��p��^F5OLL޿}x��}�7ݴ��.�F��M��^��c��>N�=]qҊ�xm�r��dV�2m�K�oБwq�H�"��YN����e���6s=��fE��G��B����TVW��j�W~���{��V�qq�ky�����*�>�/����U�<0>u����O���7�e�;�����bK�B�5?|	�'��>A�\nJ���ߵ�/���Z����1 k@-�WO��]o����h���k�oR��׼�����i9�&м�H�~��c�HV\_�ٲ��ıG�X_�C=�c����waZa���{�]��\/������i �W��E웨"=�8̒gql��b̦�e'?&�XY� �$�F�͘�ft�a�}�޶hi�aA�l�K��/g�6+J���7�+�.���dX�ҍ��+V��o4K���/��Gʤ'M��րz� ������i��>_c8����{|�'`�K���X}�
��=���C�������=A1��R������YP����2����?�v�3m���b� ��5`��P^��W��Za���5��2'��_רA���X��������X���k�e���+9��~�<�9T�w�I�Y!p%<7۫mk�@��b@�@l�:ϊ�+Μ)�
Y��d�� H\�X��,�d���b����;��P��ϕ�j3,%���:��n���"#؎ϡ�ٮvg��v��}Čz�����$A��r�����{��W%�da���9?����q����;�w�
�?|p��֮bs=�+{7\����t98���U��;_��}�	hZ�݌)�`����z�׳��<W�)>y�p���e�>EH:&'OK H���q\KhW> ���,.�l�$�Eߓ��'�#��Y���ݖ(ɷ(>@��Y
%T9��D$4���"�5RH�x_4~ܠ,q�L�� T��c��iX/?�+�}?ޱ��܏^�����Ç�@�K.ܹ��u67l�|�o�ƭ?�@��(�$��
1AM�,��UHV*��N8���,�ٴ�D�>���M�oFVrc|��<�\
WN����6T�*:�HY��
+�+u�C�Ijt6Q�`�
������!��휏BwE��\4�}]���agn�F����5��o^w�����g~u���$��w［��QM���o?�[^>�hݑhI��������$H�O��t�5�LT�Y�j�3�g�Ʋ]�܁�@/,V���x�I���D8�4C��>~�G?@�O��nQ�e.+#D�6��9 $1��׺>�\�܁b_7"�[�,3��͞�7T�{t���Ų?z������#8iC3���N޳*Wc���mcs�F���z{6�v3�\��Wi� ���B�Y�*x��S* �E�6�X�S��sj���,�)B'E�"�T@id���A�����B�o3F��	�~H}G
)Nw��^�����w����ci��p/"���v�Q��E��Gd����,��&�̺)[�Q��w�B;@.�۞G���p��g�ueL���{��U������W�ڹ��������S���8�5G
�,x�'	<�L�m @,1~RpP�ߦz�R=�PR��9$�tĎ�D�����f �:׍�{��y�E�EJ���a7CtPOC	�Z�B#	�vWP�@��m��FXm�:>-.��N|<U
���I�v�Q�CSŲxi�,�7y���%. �`�$�g��~�W�ʅg�����N�s��UD5��v��e��B�u�~��x��&�c%O{t�;��K�!F�₇�h/,<7:'��)�s��-�b�� ֖���ѿaZI$E�Ŋd'�-��f�2\$Q�Aι��mX�t�BD,��σ&HjM�&f`�h���*DN
��C�hٌ˹yZ³S�P�m���{Y�,�b��E;DOPEe�N��I�`�G��޺v�0������쵝�b�_��s���C���Ԥ	I]�m�Z/��E��NX������8���y�z��R=%֝�=4Ys-лa-j�,y�ܰ �h�6>�	�j(� ��2����3eH�x���aؚ�g$�(D6-^�U4���rܲh�"�d8l2ta8t؉ _���}���6q�y���!���vװ��*�����1��֠)�u2�I\(Y���Y�)�9��>&e��*�^��M��wX��au�.w���	�TD�r �����ӋHkM]0��%޾�w���(J6�$E!��:Z3q��ʣ/��D�b7��
B�����b�tU��f�nx̥�D��#��w/�k;'~����wm[;r���o�e���s�s�kY�\�7���_�"݄FB!���ȚY���B�b�{	>����k�+[8|Um��X�0�LB]��;��� 'G�����>:�6��C�l^��e����Z(`W�R�D'Q��qe��S�l���8�I�o����CY��#�L�/�o���ɟ.�h���)JI�I�ϟ�u�?��w�$�z���o9|��n���+w�8��n|�o�̓uX�FS�Y,6԰��d�RF&�D����<G�a�E	�ɍ�����]O���Ti�MHԬ�H6��.�j�H��0qcD���]D-Y錕��>����&��������-{7�Զ��x�7J�'&j���p"{`��Q=������>����$?��k�w��n����[����w��_�_{�%��x����b�J�lO:tfW�&� Ȱ���7���Y�f�+1���>P���)�0�
:Nd��
�����A6T>(��F��k��HWh�O�
^�ib`�]#�#���:=�Ȫb"�U�qD�)Q�=-�(�!�����U[Oŉ#��w�<>>u��#��՜v�G~q���;� t|�����&��ǡn;r��n*�2z��kzV�ȭ���/�V�+1��B�*yK뿛�sÕʖ���zv�	tl����>ك�
��Y-�?��}��_�����\�9�$)|�ȳN��v��5O���]���z�U��������    IDAT�⤑n,��'n�:2�/�	+�������;��vp�<P����p�xj�qh8� �1�7-)c%Q1���-E�x���6f�i��w����u1?0E����uo��b�I�Z� �c��O^V�)��.EJ54]!d�?+Nॎ$R�^��KÌ����
Ct#�@PC��c���S���nԀ��&�n>wx��E��~��#>���{z|K������ _w]�6�$d�.�]X#�G.C���tt���8>F�!�(���O�7�����ݴ6R��h2�1��yi�4?|����/�,�T��Z�P<+j��`ua��bqe�$�X��0��z��~�՛��R����9���]d''�O�t��������/�E>�h��q�dj�	�I���nZ<���	I��@�Q�5���2��aE����ܡP����%R%��_���>���d����L�P�ҍ���V[�q�@�u �؟�ŕ%���C���6��#��^�Ԓ݈1�\D�ԣ��������G�&n�>:��U��v���p�<P��!�����YLS�$�r�K?c����fҴ�@1J�$�r7iVc��~�b���(�t"t�(�bʱe3U˓��k���=�+�d�|N��rl�$_��6�՚���V�(��f%9�Rօ%�_z�^�l��o�XIr߲_%�A����g�3O�)k���z���W���xU�_�{����-U�=����5� �^_�ĹY%J8l*Ptd�*���D�DYc������rᔑ
�[�*z(�!a�Bt�!|�|�m��u `<� Q(�<M�;@�GGo�l�� ����L1jSs���4�t�i互����|���e3H0+*s[+f���X\@��\}��q��ARc��_�����3��e��]����E����wrq	x��x�P�樋x��h���RY�%gR���@.���4����C�� �����_	M��-Ӌl�&b�� �t1�<�֍Jx��|�d-m�P��J6Sf�|�-��.���`�<���dE��=�ԕ��3E7�7Ʃ8y��j����Α�/��}�
���;ǼE,��s;%�$ʖ6����$��\�s�I�
��,Ԑ�ug87 ��k!;YҌ�A���<�F������n��t3���f��!�bI����v���)X�fP�s��[�]����Nqq�в�1�Z�
�W��H�1z�D,^=} {�� NY/j�C��M^�ct��1�W>��X|<�d�X�%���U�-*�;��
��8E�|�|C�W��4Q��h3����1J�� >ގ�EZm�51�E�Y�I�Ǳ�մK��m���������i);�͉�4���h���2:*e!�h�"5\��1RZ*����R\�>���s� i჏�M\�}t���[�����D-:Rкs���M0!�YoU�������Q����G�4����1�/le�B�e�Hb�����X94b��J8r��iz����D6�B�l�>>;�P��g�Q���Z.�BH��"�$J��)CYmT���@����b��W����:6q�g8y��]t5[-Th񙫩s[��4����$5XCd�Kȭ0��Ol��g�V[�BNA�{	 u�9F����̧��r�pҚ���x)~S�`Œ�;�B$�s���ag$T���B�j� �Խ��6#�cj�+�3��T�?���q�T����ˀϢ�n�o|V���Q��fk��H0R6��B���%Jј_DTgG�K
��9u(�͵<4 =����WH�պl�$�\�ED��%;�~[K,�sp �����-DY�l�=>%���@�z�}K,���1�lfՊ�\��,���NIb,~���q�H�����&�^�ş}�MG^���{;=��E��7>�!��3#(ԭ�i\f{����T��)�^R�c��[P�<������ۭT�#N�P�AS?�j�α`y6�ŀ��D���a�"	#�T4�(�3���	r��{���sm���5Ց�Y���iT�Q�4�0�쏱�L��>6��=:1{��������]�Wq�i�dq�ʨFbw�0-���,%OK
[M(I��@s`�(&�}����2%q(t�"�6�왢��a'Ķe g�!	5Cfe{;����24�oR�"/'m4�j|O2ef�2<b)\4��cܩDR�5�V֫RU�`=����~���tb��U鎋�+x*�.E5��иg�0���o7V��Igx���$�gmEm3)�� �8���T�<���ֵ����������|��0^�6uM����\]���i�Z��ո�
��jJ�+�
C��'p���;����L>26�g����[��_ݻ��w�����	�Ք=��8���◖�ѿK��p�z����l/�$5|`Z.�9����J�)D���uǌF>�+2��~��{�k�R�G��i�[�.��׬�����1���F]A����j���|6E෍�"�7�W<���	��8��K��I8��N#�/n����g�3��MX��h�S�NE�u�S�j1��GhZi��?S>3�yaV5Z���l�	훹�xC��{h8��Kd�
A+�m�ŋ����j�щ�+�[��?��۶|n��{;}{}�Eמ>/��Ǟ�,�� F�qS[v�w����/��u�P�Bb&�&�⏳
�Q�1�1��)H�i	���%cu�T7��0�Ȍ}����BWcH���3�Fh���7Y��\���z�������-��~������ڪ��+|�((:�����V�c}]a��G�T%;d�#�g�	*3ф�ˮ�����uEIJ��wO���;����C�[jy����/�%	?'[!1'K��e��+�'BSih�n�V��l�V�2��W��͵�>~��Wn_�������8����'�E�O�Wg�MǠ���'s�x�O�9f���@֏V�b�ו��H,[��>Q� �2 �(���]y(�ߣT�P������h��☠�4�k��l�͗-�Q�4�hUZ�u!C|�g�D��NFB|-z�h.�c���R�L#t!�P��g���m�){�����䗶���!�_�؎{���,t]���q��=�A�$���̠\��<R���\o�$'a�FZ[�P���m�m��R�$ś�"
]���r\��X�V�l�'��:svcw��9�/q<+\"��R���'�����+���{
�*!�ӵ���(Z�g��}�^�M)�Ӓ[��^a�UC������>��F�0�0����U��>c����������6*_���������Z=@7�VΊ�@/��N��v�=�w��i.}z�b~|��᧤�Y�O$	�+y{��%�����AZ���/e%Q��������7�k��IZ+@clF�E�u��"JO��pz�(�t!a���(*��s��-ʥ;4��k�}��9
�4@k]����NZ׃y����_{��UB��?���N��XwP��;���g�nX
�Ć�2����1�!"�|_~gI��f�"�%X�B��D��i��vl�@g��}��ss����F��,�V9(4�t�M�j��.#?ЭUk�n8A���H�8GL7~�a�.���N{���!Ǝ�Q����� /
�27��z�d"A%��ZDy�W��������O<66��sF?�2�X
i�����en���ڛ�J�|�y������K�2����Í�$U�a�Aa�N����i-��E>T��O#��9�Z�ck}K�p5ý�$HI��[�j�uE�^65��<��"��%{�x|�4��%R��ؔ�EL�d�NH�a�{���v�p��m,O��Ccb�̢ɶM9Ѐ#�s��BE��k/�0�K\}��8qc/��ӏ�OmU�n���vz�Ɩ���}{�G4�-^�6�jM{�J��A�An�KX�v�`�#���)�����9��X�P�ޥ�a%�<ԣ-WƩ�(q
G#�«�@3@���f�:*5�*���ݢ��)�|�����D��4��	5!��DF@�I��u"�ۉ�����$�c�H���6�t������V��*�c���&���zh�������>�R�x��Pw��a����bRC�-u1\�:�U�O�m䆺E�(�8����V�o�µr�Or�"-^�j�����Z+-�>1UQ�J��rv�k�ʹ�=e䇴��y�2K��� /�f��Y�7���N������B�Q��;F��Gs|�|���6y�d̺c�Nw���5�_����M}Ҋ�������չ���dc}�F���{��8�ht�r�AҊ�劑��j<�8x�"@�j�$�I�)�H�%K�_�R�;���픕�q�R:�b7`/SS@N1�ԙ-��j��Q)����q+�0QJ�)@�O����4�E������]�&z"%�8i�	8W*d��a���I"����k?×.<M|�"���霑�?]�';l�]����^�]?��Z�E
�H
����L���5�*o$�m�\����5�tiDՖP�I�x�j��MBQ��;�hš̕��ؔ�?l0P��J��`W�X8��q��8����xh/6�#�ь�y�br���7g�8훕�8A'�֛p)Z5Ml:�[�����=�Y�i_��8qTz�f{m��s׍��3s���m������[��9|s,B����HK�N=�}�zɪQ�Ғ�dE!d�+�X����;�������]n�t��04�����O�IXb����L]F�e?����(�!.ǿPR�H,e��!F�V%�w|�/�-mAzs�����^�B_mͧ�%g�>޹a@[�����ڶ�����U>�o
�m9A���ڢCaәvY�e��tI�h�aM8�x�T0�+G�HN bU��`}n���K�=Z���	��AϏ�	���T�d���c�l������ul����Ϧ�C6]~�XB*�C�N��]��y��Ws��㔵}h 3M�p������8�s;��+{��E�������6/QJ�ڲ!��4Ѥcnޮt^H��ٕ̍ƒh鸘��O���ZFk/�Ej�Jt�L�u��
��|�">�F��}K!��Q���\��@� r�2�ȬHC*���D��bn�RVc�����q�_Ӈ:0���&o8s��Ớ�o����޾�h[��ڇ_Ľ���o9�4F�腝8�H�7��W K��X�������S�hj���d䕰�S'�2���=��N:e���X
&�43yI:�djǲ��B��e����F�*�� �C&4^�L�$�a���Z}60���_r��;G���_����uC�/Z=�k{��������.Z��G/������v#�+�{��>�X�гe��Xe@�&פ^k�dE�kf���QF��$մ{�>����\����(F���/i�y�\��ܢ{4��BC��^?��^gYe�e�]��P�\�h2�dm�O��3�#�1"��CO���쵫�
��ޗ�ZSs���z	w���	�!����{���ŋ��]u��$�**A�*}#��T�S����Pe\��"�L�XZ|V����5S����T�$�1�����9"��͕�,�5+�bW�� i@�G�BE��l�By/���*�Twv&1�Ϟ���o_�K��'M�ݺv��)������-������i�G	��K�q�[_R�I�d�ܬŝJ2��nK<M��F=�L�)�R��9��y���R�M�>ڵ6D����b�-�Gn1�)^^G1���ސ�pn���[Z܇�>�l���Z����5�u��j�����)Y�/������vM��/��A�c� ^9���m�׏~Z�����-�b�"����������_y�D�G�m2�fhRi��Ġ�d�pF�:����S;D{v��	�<�v�<O�����D�RB[�����3 ��I�����!m���!��i��Fs~QTk��ٙ��h.ɚ��{�WJ��$�O���|1��ZP��|q�Y����Ta0i����p�Eg���Rs=t�����9|ʀ����V,�(~�{/�g_A<�	��1�+$n	���1s�V�.��>�*h���OL��1x�F3�D�>�"S�k��(�Q��;��e#q��a�#,��@�#<_\�k�M��T��~&3��3	�54g���A�=�?Dv����׉�@/���z��Xh�,J�&�>Q�qU�f6�F��J�Y�����>zNڤk���Mݺut��ǘ3��x��}�
]_��K����G0����K���W�0�-�����
6�C}�*��u乙�/��� }QvQ��`]F9��pPЇ`񀀒��iEX84%}�yΣ��f3��p{J(q����C�̦�܄`��ִ�H5d�����WP���7u8-��h��К^��h�hf��-� G�$��Zs��[|��g�#z���<pp궭kW�Gn�m�%�ο��Ɔ�E�W��E���kB�ʕ�ZO�3�G��ʮ�������Qh��ԒuNӈ[2%C�����դ��?ܧ���C�%��Q�5���0,���>��6�������/�fƇL޿55/a���4�m#P1��P(aߌCC��i�.�=� ��S�lJ�BqH��J�bE(5��1�K\������d!d|j�y��h>#���qw�go
t寞�m/D8�A/T�I����\�v�5s��N�@��L�&�w$��3j�@^2@F.2q��/��ŋ��|<��z��伴�ӚɩH�P�a1j]t���G��n�/6dop#����ȩe��`7��w���'Kf��P�>��d���_�-�ZH���Ic�U���J���W?~6޲�"�?~h��UY<�����yO�����|����hs�0{L��19��
�� zr�}ȕK�	ډ$�,rj���tK��� �y�sC��=4�3	��ޞ�JD$��l�^�C���k�Dg�=C�7SsYk!�Y�j�8}<vˊ��v*}}��8&��؎����ٚ�$G$�&�z��4�� ��sl������������n[��9s�]�?��}�9��l��=����-ű#��f�����5M�L��%� �"�3���:�`��Xg��jn���A���Sѕ$�@�1#�v��ڄ
4�#����]��͵��A���b��Q*�y�X��H	��->�p��.
��>ZNֱ�� ��jSJ�z�$�Ճ{�J��ʍYx���/_p޺����GN�ݱv��7W�y[���[�@���y>ր��4���VD	�댏7D����,,p"�4�AZ�!]VI�o��Q���'R�Y�tx�g��2���=b,�SM�0��;�A3�H���e��d_�bY�o�\W||ģ����f
���7f>`��Y.̨.�^O��
��P?{
{���������uU��}�G~n���{}�ȹ�_�����t$$�b�2������K��m��T���:nSgi�&�H\O��RN͊
�+O��4%2�A�]�}@ IL	�cE���8n��%��s>�]\->kl�7D#�M<ʔ](����G���Y��@��s-�����ܴ�A��C�l��	$/>�=[ߏ��t���m�j΁:��[����t�]M�5?|������(F�+��H\�HR�F�(15/VF���J��5i�!��e��LL�bUZ>0� �����-�,T3f�J���KIR+�tƩ����b�jgC�c+�^#��L�'E(3e�����r�B/b�6���$�8�x�h�t�=>6u������8���o���Gp���<����p�=	)��h��1�k
�5�oTs�:͖��pLݙ�&*r87�	�Q�F�ט�25C�q�g6{@,�T��F`'�i� �yF���	=�HOo��)&f�/i��CX٦/4�����C�b�����'�3ߋw��㏏Mݱj�?u���=�{g_��32��9�D�sr���Á�8a��4���Zy�{�h`����7A��+1�(�+Z-��8de���P$Q�)lp��^���t���g����Z���%1��V���F��������z��~P|�)�P/��;)��cw�7:|�C$�� E@����X�ۨ1A��    IDAT�?�}��Ǽ�5E��w��Q�Ƨ�5YJ�t�-���V{fP밺֭3`r��'����0�l�����z���z��̣ٷ�53�eQ���
��Q�1�r�b�������Rd5W���gGHsx�'���i	���غv������z��>o��n�=���������D��Mq3ƅ�0����u��ɨG�9R��2�$'v�Ez�^��MOl����'���������׭?
:rR���x���7K=w&��.S�RN?f4#*8�B�"����������lf�ѫ�5�a���'��p4֡�cwl]�ݺ��ޜ��ʞ�½�xo!�� �!��_1��W���.�I|�X"�M��l�%� ��1�(��S���C�$��A�.ܺ�8��Ӄݤĕϡ̣�I�%��*�M�5a�,�W�h�6] ϭ�("_d�g�i���_�kė��T�Li�H0��2�+�x�1�-�?v����;��ͳ��_�u��}���f��灧5�Ǿs�fq��%e��:� �K�3fz��yչ*���VSB�45#�s��ýb���%$����B�#n[�����!�%��T����g�ϼ�{J}����:ߗZ��&U$)�1�ӉR��2f(kIh�C�:4�%�<RZc��z������p����n���\e^�.|�B��Wc��(-��p�����g]��C���6A*'xp6dBz7�J��Q�Vg�!�d�g�jI�y��j$�䙬�{$J"X���(�fȜK���*Z��I��)�!H��8}�{�$g ���X���b����4=,��#
�R�x����ʏ�fZ��c�n۶f��|C����_���[�.JW��)|}6 ��d^��=Kݔ?�w)��<��ȷ}Ǔi������ؘ�$iZr��#�Z#j�����b�&���	|��$�V�Ǘ�"�sm�Wu��F�|A�9{��2wrzQ��M���L5'��[F��S�=Q:ˉ?z,W��u�i�ᬠ�e�1bի�՜�>�����ܻ}d�n~��{;s��U��x
ߘ	d
_��� �,e��r�J�T��� 7�8E���q
�Z��d�(!�(��K>:Ga��t$�T��|��	�N�9��1=%&P�;P퓬�]#��1�$Opp'JsW�d�B�~
����<i�캗����f�\\�fN	��~���I�B�	�;V��w�oų6�l�/[|ݲ
��if������c`k$� ɔRG&�R������z@2)�2��9< ���$"
���gF3���tA
�&Y�%���a��9Nu�Ke�ų�A4^%y!�AK���NoY��Xd9U"//C�l��]��,ɒ�|%S��w ��ӷ6W-T�|�h�tf���S�T�l�]¡��֣0�����_0���	P̣<�#�V�^'���̢�Ce �V�8r�)ؕ�����\����$�U�W#S;HO8Yz��C\�O��/SV�Tjo�	c�h�`��(����o��M�=o��Μ��� σ�Ǌ,Oē�uŔ#ҳ<�C:���)�$����q��2[�uP���8�\J��q3]<�c7@��/*_�B>0�*��4�����S�$�0}��3���'��$K6���Pr	�ZX
���� ?����-�r5���R��!�Bf̝�2�i��2}��i�����@١�Z#�׌����TRI���J�ТjRO?e�Z��ze��ͬ�U�_�7R��g�S;��p��,ɓ�t�/����XvH~�дZϙd��>g���f�+->^�`2���2IP9+��+C�iخ/C"|j�I�����HL�͛ʁ��3X*��'�-5�|d*c��27U"ې^&�֌�j\Q7�(�7�)X�D�l��?�G�߲s�ȧ;�̀��Α5]o�jh��\ �e��:P5�:.u�j��3=�G�ѥ��GipR+�vMel`fE�cR�a����A�L�1 ����#[�<�㈄!������4��G5݌<`Z����3��s2���ow5b����X3r��I���l�?�f����7gåp����&�Y�V/]��yf���?IT��v���y���3y���e���\9��<O<p��ʨ^s0�t�� ���6���s��j��ތ�s���Ui�&]�K��`��fh	�t.m�+�͢��:�߱�^����׏0�_S���$j�D�����M�k��VL� �<o6!�q4k���-����.�PH����(=1*sUzh�-�c֛FRc�Q�f�p6�X�߫ ������`����߲*�'�۹�.m��of�[��Zrh�Ɲ�%Ç5�eN��6�؛dBM5�%-�Ŋ)�����
d�+�%��˔m��D���5��fX�N_��M\8xv���oK�#p+&uh���R�jVZ�
�=|h���׌>e����f�3s]�����Ȉ��Rms�O�Փ���*���H�2��Jx�<:��X�*�!\��ǰP�]��'���\9����n��t���53�X�}�,�O��(���ȯ$`��*_�q<i��?:>y뎑�������Q���F�_	<3ו�1�V����&�	Y���R���������qI��<8傜�%P1CJ��8Ak�
�}L�3k��Iauw����,.�}FJR'�)����M�t9�\g�<b���vz�g	�YT"!��ue���ܶc5��js}#�Q�-B� z��ށ	<���\۳5�g�!'IY��v`���'x��s:|9�+��n�-�9=4ڰ�-�Б�0�&��ۅ�`�h�i�d0yP�"�N��#�2�\�M	9n_8eD���<�F�Qo�9	��3��m��**Pr���m��r��լ�3�`E�#GXh7�²���ch�YP��*�S��E�*�F�Ɂ�By���qp����#�O���ɢ�!���sJZ$׺�Ҙ,+�U+�E���x��J�8,N�n��EGWE���]dr�7{ ����j޾�W��=2>yێ��ï@m�����Z�w7��\�ç��3!,��`�h3ő�lv��f�1|#*	({a�+u*��l��c9//�8E����e,�w�+���M�"vu�k�"n�B�	�6��2*����@櫨M�ie23VV������C����:�Ǫ̇�7,Mr^�Ö]Mo�`�6��'q9iᵢ&ep���?}���߶��>�;�t_K]�d��'bAx�D��hy��4,��kI�P��FN�4�x�a�4'n��>�'U��̥�^���&7��l�W�H�¤����KB�O/�*��G�%e��&�x�U��ѕc�zB��V����G����<�k����2P�s��Rע�H��'	F��H�>��v�N)I8��j����7n�d��{z=)v���ib��o�3��㚉������yt�Cc({���-7^Hlx����N
��V�{j�la��Dy[T\-҈�e�s���A��43v��G��"���&ȸ��fP���'/CFYO�� �p/
��,�K���˾^��6{��MR�	F?�8���a7Zfc���Swl\�v��o���]�����#�@ߞ��}�u���DN	�h%�/��)�
��3>�����.N4'��Z�.�$�N?;��3��I%))�w�j:��U�ˆH�s����͜ʴ�$�%�9W��㊣�O�k{��	�w��S�)���B��f�k�NF�='�$�_��_%X�XE��Gqն��
�H�?>5u���U4&�O���N��\����s�7YA��0��Q��m�Y�+S���Ŝ=�I���@��c-4G%�`K>��Cȯ��1��X7-����y]�ʕ��	4��S?���?�b%�)����!�BN�z������m8C��˼K9lQϢ������2>Q�;���º�*�>���~o��p��O��y�p��Y\����_r&���v�ѕw��{�|�9쟬��fQsmX��9vC�c(�x���*��/&�x%�[�j��Ko*��8�xo�G&<	ݛ*}
f-D01/.�S�-���V)|=뇤�A�^I"��8��-S����O�M���@����1Cp�(]-�N+֓;2Ά(Tmi0^S�"�ɣ�f�ix�@Y�?pp�έkW�g���n�,�==�{&�p�;�"�%��w~�'H�nx�VvdH�M��9=�v����6�16+� ��"ܡn���h�D?0� �X�e�����w@�U]���U�չխ B$!	0�`26"YHx�a���x<�6�q��	6 � !��Q�PB"�b�s��ʯ^���?�j	{��㿖ׯ�X�T�]}޽瞻�>{�tyF���y�˩F�:D��Nr�f'9S#����,W�����PKr�yȂF��2��]c/WP\��$( 4�k�X�1"2s�v<6�˘X�+�}{kǒ��${f����6kY�W����������$�v4s��q�D��p0�:��ˀ,�d|�x5�8K`��	3� �x�)/b�
.Ei"�R�DR�`l'Ln�&�$�r�:����/�hI��I1�i�T��F�	J@a��0�">���3`���)J����8��H�E�ܳ���
&V��Y�����3j*>wri��6si�*��I(x�]X�2��g"I����]z��ʌ�e�� 
ޤ��?j�Q~M[��Gy*D5�'�)���'�jZS�IG��t�sM"�fn���#��3$�%���r�H�L����#WVӨ<�ϣ 	)݆^�?�c�����>w�N�'�q}G%�-!��Bǉ�ٻ�Ι��k��j[s��[k*>�D��K�!����'~��nzfI��dkެ���X�rV.T@��-+sIGWw���ұ\X��KKW!�ίs3���YA��c�E�$�����Ii�{�!?4jZ�amf��$0�I����x��&@��P��Z繬�OH�A'l![)A7�ZO`�9�y��5�Q����Z�W̬����Wř9ci�-��5��r�f���[���
�")�!���w���4N��s�/�:	�"~�Ԗoa�m��a6�.X��:�{$ʟ�	Wz�B��"�¶��Y-�Zz/�1Dڇ�� p�._�U�^<h�)��K~��b�� �6~�qZ]!��;��t��Y]6|?W����[oYZ*)c�r�Z�6~�n�j��u�̦�x*�iYŎl9;��
Hd���u��f�"u�y�2yi��-�I�b'����Iu�	r�D�{�8��O�5vd)��
"��پ q賯l����#pO�_�Ka�A���އ��<
|��_Q4|�k.l|���ʡ����yz�f�b�F$��@��HdQ7�_���]Ek朻jLپ��z��/��mb��#3|)rU8�$���0g� f���-K��z?�F#{"�h	�?f�閻���hq?i���!89{n��;�r.p��9,9��y�@U��S߽�GV��v{ϲ�V�<4�TC���;��:�U�3﹭��o!&���H��!��?�O�&��R�Q:���`(�xX�iu�<:�/�"�C&�Tb�3�q��Oe�@q;��<����yv�)/��.���=լ^~����%��߀��q%k�� j�$<���YSH9~`{W���
��������V�;��O�~~��Ĥ���*�*��B]3\ΞYr��O�D�E*e� �
���`��>T��E����,�E��W��k�P%�N�H�Y-�5,��� ��?64.��N){���N�d�NN��(��m�5Mώ �CCr�T�Kx�{�������n�Z�������sG��mw=Wfˣ|^��]�?_�Qx��y)������^H\1���e���R� g8�:RLbO�,?]����$�L�� F�������Hw�A4C�� z�a�FI����%QZx�q����^��L��C \���,?'�S[��\�w��R�F��t?��<�_��jKib�WWx�W��v�����G���٫K,�Q�T���7��5��|½���O��b�إ3gm|X20S��%�{hQ��!n�ODX�?$�L*����JKP3���D�,ĉ�	?�{����i����Z��I����8�d�@9���?vB6I�	��hȍ^Cw�<β�K�u/���T�Fm��|�A4TM;L+�������������XU�(�UE�翰?]�{$=!Hf���t��H�&cC ���u7 !7���0T ���\sl�"�1U6�`j4�M�i�0/��@
�
&����R1�}(--A(' �����b14wv�?���菥q��GOt"�r�jA~ L�➁�ϒ��鄡 7J��h��4�t��� I#�v���l^�f��QW��3߿�E���vv.���|���v�����UE�:FQ$���U�����c�gA��f�, )�0�U��4����Gj�d�]�`�8�&��Ȳȿ�@~@��3ǢЯ G�QY^��'���|ι:Ԩ��m����׏�{�E[�� {?8�ma$Ӥ��3/4�Xǵ�&�%�.t��[�ĔJI��,�ȰL�11�,��Дx4��b]�xa����(/��+������;���U��E/lÓ+_����x�F9�](0�5�B�%qYB�ׇ��<t��a�%�[�X<�ϛ��Et�q���2���tz&�>�è��|�8��~n$�M�N�;���M��{��{ch����v�@�x��+QA��!3�S���D��ꚼ�����~�8�H\���0M>����O��cь#>G��ٳ~v����i�c��xv�+ȱ%Tv�*ڃ�x�P�a� ݤ�����{9�8�W��P%bz�h^dIL�/.jn�!
��(j�`�x�d4֔b��1�,̓a���u/�`�M9(�;��J����m�[���f���q�H"��)=:��tD��>�K�?f�={�8�Hi�C5�3�:��Y!�\�ӊ�?�?��Њ��پ���ϓjN�ٜۗ�KR	X�\�K������q=�=Ёq�>� IiV�&�
?SR��	�=!�˯���Z��
a(�/�f�9{t����6d3�Ig4b|c�j�\v*�sY���,�I�3bt^�[��`�e�&�c�G��x��"�����&�&:1�S�h�	�D��ŋ��{ 9$����L�3nCx��Dc)V���p����پ�s��g�=立�9?O�F�}���c���hL�0��8��kECj 9�AnT�⡚���Я�q4P�=�#��t$�!��a:��E� ������W=�;�+/��␂Q����Ӑ��no�4�U5ֆ����+J�����$~��F�ŀ}����N�HG�E$ĭW�O^���s�5H�e^��%M�O�� н9��p3><�L����?����g�W?�_;w����k�ܐ���
e���X�hΈ�qi�A��ߎ�L~;��R��YhX�kqME����x��U�;����'MSQt�9�b��Pٙ����z���@��d�xL8��Dg�&A��x�\�a��4b�q�B�@,�7����(>n����à��V��v����vX��d�H#�x����P����~�^��a&|��v'V�}&�t�:%�^>\�x�,���}Ѭ�ϑj�{f��?���gr-��5�kV���<��#\~�C��o��I��:b5��KhR�T`P+�o	^)�wK�ЙW���fP]-�9h2�C9�J�(j�sq����X1\��I�xZ#�t��uHt�y Cu�>(�4J����������i�~|p��=1l��.l-���G��� �'g2,	�Q��O�#�P��ƫ��`$S��<�{�v�{���<*��gSW5uǶ��.�YQ5���%>r��ge���r/�|�-X�I�(~T_;Hq�roV[�\Ro�V�w��x�����Š�f�(X]$1k&��d^�Dy�_�6���3q��1 ���ܥi1f�.N���+�A��'MQ�mڎ#h�b��}�h�2
dO��P�,E%aI| ��|:��4t)��E�IB�t�,i9�Z���c�DQ%؉(��O?�Gt�    IDAT� j��nlm]2����_N>3���̹sA>�Hiq�so�Յ/��X�5DCov���R�ˁ�`8@B��R�(�e����
�� ���j�i�� :�J��l�zm\2m<
��M�)N���y�5'4U�$	E%!�/Cz0�h^d���o�XO��b�G`�A�,��asS��8�S�۬��;�E�S!_���h;<��jM' �[
'XS	1��W�������o_��`}��[��.}	c)��r�{ZP�D �C�au釈���V���Jl(n���r�zu$\su��m��,��R�0rt�H���btu1�su\s��5����	Tt��B�\V\sL 9+E��M����>�G��}�8�tÔ���[��BmK6Guab���tt�� -�;�
��NY
�z	2�Z�J65�5V<��/~���O�fc[˒ٕ��{�_��S��;�9M����s�ְ֡0�����aL���Iŉ�r��]�������Q��r����'BE|���q|�T�k���t*�j�{�L7ZzW_z!�H�����!����M���T*	�W����ځ�[{�Ic���#�D�R�j~�*x�͵� �)K��bHx�t��`�� Ci��֋a����C|�h4&�
<��> ���e��
���Y2��w�^R �":��6a�җQ`J���i��83܋�X/�f�er�"-+�u`_A9�����*��9B �	CbCu4�z�Y5�I��N�������DYHCCu	Ι0#Ja$|��<�	�'V �yTѐs�$���Mغ��32�i�{G[�5D�!G�BB�F�41�νlJvȎ"������˰tJ��
��̫�����@�I��uj�7��,�U]��a�x
��@��jY�f3�Z�;ƗƣhH�1n���A�Qx��##%�мh
����ǂ%��KS��� � �1~
����FZ6�/�Q?"M��[~Lm&�5^�
��_�7G���y������v�F�ᠹ7��?<���ٛ�(7���5W�&��x�r�7T���t?�p�t/+H%e��"$rj���L�&E����w��H������_v��[8���}y�z��Ek���I��tefU�k��	xYt�h�!!i���pܟ�^_>�RH]@vR�AN�$��Z�p�0»3P3)�0RM\8y<
�2�|*�F��zF�(g�$��m�kWW:��GN`0e#j�غ�#4��T�L�r���rH�"K֒��x��~@�c�Q �����oR�!�+D<T��L[����œ��u4��e��~��i?���!u��ي�V����f�tL�)�2)䲥)�*0m��I�**�t?R�|"�߸��xw��!%k˄��iґ �A�����2�	v:���
��A��T���!�!K"e,����Pk/L=�hFB�v��2m��7WS4g+��(�sI̘���x�B� ̾f��n����ǇLN��#��r`�m�h>6C]���^|?���ںtfU�=�^�7�]p��d��L[��V<�j=%�d��L��qy�#�� ��Ml�Q�Zu��Kj6C�{<O�������בJ%�htm���v*|��=�p��F�"���@!7{�O����{��ЗT1H�O��H�ܣ�L��V�V����(=�\2Z� Cjt��m��6��Nԕh�:�'?�� �b:,5��P�8�� �
�x⻔j�H,/���}�5����;�,͵QO���/lœ��#I+���s�͌ߡj�0��*�V2	�y`$�s����	�6��͈�i�bcUm�w�P?�#hvRr >���($�M�ǫ�.==���6��u!�p0��`*�?��4��hE	h*= i"D�>���S�-�Ũ�qh�P����T?��T|�(͕a��;:��>��>@,M��*tՆ�x����G��S��-�Kg֌�����\#)�K^܆'V�q2�y�=�3��b�@�S��F���u�K�Pa�t�Ɏ���5B�t�2c޲e`DQt+�pO��/��P5����\w#�<t$2*�DR�u���N���HkG�Lһ��K%��cC�����"W6�� �>f&I��k������6�iA:�2������7��v-�QUv���3����]wR��Ʋ����r&bfU�!��CY�Y�B"C @�n���"5=����J[;/'�d2ɿ8�Sx�k,v����SL	$#Q\r�6 �>H�w��#9�03�Zl��~Ժ��Z/g`gҢ�N�^6�@�鄤Cl$����A;��ݜT�ZS&4����Γ@k���	��tl���i����v-�KO�������C+�(���D�rLa>�Y,�ܽ�D��u]p^H����h���s�į�m�Lb�)�qH���ҧ�h��D<ʔjI�7��*��F%j:%R��P�'��OR��N������g�2ԧ�0��F�ݩ"E��ݦ��u���I�>Ē�WBZ*d)w��h���xŋ�W�~�@�����`�~�Gs�X�砖�x6
g�����cW/��Q1��tjJ��;�pn�I�]��6��F� �o,И`s%c%#�T~��4�Y���x<Ν��N2���Q��dS��~`q��i\ɨ� �	�^��!�d*��>=J3�V���a>هB艫���4��f�t��_�*P���O�)��� �p�ڍ[EԡO�Eè����c�2ץ���4�e&Q��#�̓p$���5C���Q���9gO@,҇�`���Q]?�7������Aa~���w�ť�z<�����i�2��-�be��َ�����CQq���}�vs��o�G8�#ǚ�D����S2���+�W�z��7X�=�ë�E��p�OW�O;\ͭ-�Ko]������'�>ˊ����<r�]��)��w�����J�����b�����È%�}�Ty9A�8�zx=�g/Ǝ>��8om|娭�B2a �4�t��H;z��}�fނX7"�}ظq#�:k6��),_�N=�_s!֭{�w�ă}�T���_@�������[nB*����o��o���}۶�@sk&N��@n�ܴ��eMy�@����y~2�5���j�F�X�	�'���H5�r��WkKKǢ���ð�����9�dTS�����d\�
H�&�Hg���1'�T�PԄ���lg������֬aRR�2�3�\�;p >Z���W_}�]w#v�އ��?�gt�h|���xq������_(���1�ՓOB��{�]���U�5�1�v�����w����������)8}T�a��#/7����U�V��ӯǄ���3� bX��5+����W��� �B�b��.l�{���w/��R|����֮�3�?=��O����Ͼma���(*�b
�U\��>Ç�L=Kr���睃�ϙ�m�7���f���c�%�}ƙ�{�9�}��Ť��������͋����k�c�z|��)����(�^^�t4��������K/ƥ�_����!۱�}���z���$)�a�WoBCm-�y�i\u�u8|�0�-^��L��Q��a��u����@,�j�P�I!�sr��;S%%T�L��	�:������v-�u����]�����=\)��̾mQ�X�x*�<>�:��3�>Ьt!��뮺Ey��{������'P6b


�C��{���7�'���Q���ע���D�w��eo}�����|�MX0�)\~ť���EM�������{�{:0�1y�d|�?��s/��\rڎ¾��a���9
�7��ۻ���q�fÛ�F��r�8�d{�T`zJ �AZ	������j��TC����=�N5�%��yЊgr+�f+���̈́�H�0��'����M�p����M\��]`N��#5�[T����KO}�h0�J0�E�j��De%�hm:�ښj�w���dYE-�Z���}H%�P�4��
�����	[�PQQ����G>���q:"ho�nkJ�� �d7��m�ak��x�`zk _� 9�RNr��̖֮E�+�7�[p�o���ϭx��&l\B�k�N;9A�+_�a^Aj@��{�|<@�1�ׂ��|�+��@�t�l$8�v��*(2D��.���"ܪ�E�
�w���&O�����ؖ���d<·h�`L���MAaa>"�8��$<�|H�FgW2
��9��3��������	Ԡ?��O~�:�o�,�g�u�xJ5U*�d�&���t�/�y:6@|0�����X|� 'F2A<��N}4�d"��B����"G��N:�&�T��-���f�1]CV��_K������2�7H��������#�����������M	����4mA�����ԅ'%��2�JF#i��4ɥ�C��)+� ��3�ʆ�N~���o�.ٓ31rM(Dͤ��tF70�'�ʸ�$�(��t<��e���%(��GNA!�f
��툷q1���S!k3A�<Yj���ha�*��/A<Cg3��!\�8����%B����y��r�QS݈|Ұ1�v��� �D�&_2z)d!j�O��Y���kѭ�e�o�p��PB%��lU��(HB��Zw��2L��'X�H�)t?�X�	H�$�� <�X�NB&ȁ�0�fR�$	��=:$_������ 2	�?�N J?'I��3���S> ��Q��I&�}���g�d\v�y4^ȁ��3Ja;2�`!F66"?Ǉ��N�d�!e�P�*!��qU���� 7BNY�m�gT��;|�lނK~p�틋$��|�V�j%��~W@��I4oJ��P���,(�+܅�����<Y�@�,f�L�`ኪä��B�н�B���'��8m�����T$�%i� ^�r4���fRe`�C�Ʀ�(�Dɖ3�%D@�F��kG���=�'�d?s��	"�-�Z~b/�f�&��0j���bj��6�t.�U]>|�U5?�m֒I��մ�|B�&��(�8Xq�y�{���@���a���8ĎC̂_.S�Cq�@�K1y��Nz�0���n���	����C��l�&%���ÌjP�7���׋�^.q�����#���2� ^BFA��PUƞ>������BF�q�7��L.�2����
|C�����3�J�Oh��Ϟ��@��p����?I]�f	}0�VP�9&�pZ�o;�e�Qm���(�w
�2����3��{)�f	�1�:H%8���q�~�4u�z�����*OsӥN"�u��mO�'6Қ'man���G:
Fc��s���Js�+C�`�+���������@�����T�������g�j��5�����G�48M�9$a�����(������NI8���{o��r��uUE��"������)n�I�άf��@T:D�3oY={�q��8m*s�mL�x�`��Q��yzĖ<ȯ��'N�7��M5�D>^߾+���_ ����TC+����{�����3�̞��@���J+��o��u( �́w؃�h���D7d+	6j�UL����J�[��-��\3^�Gs8��p��Q���X&i�U�$!�H��&ġ;�%q\�W��@ ��_�������P%��L���c&NC~a!<4fG�������D�bf�l���H6�<|����/	��f�ZT,���pݎ_����B%�<�e�^�m��q���eF�д�u �]�����L[8}�xL�4	�dc��{���}ba�"�.���`�m����S��������~�m=tX��ш�a��DEPV]W��;yyk^\~���B��l޸	m�\�g��;����h�0݃Q�|��%1��E	�r<�B�W�a:Y������Ɩ��3�?GUs㼅���;�����K��'�L���j �@O
�h��fo �<�k�˖p�]��o�{_�^|�9<��\�~� UلO���(Ws�RQTR�o��8w��H&Sx��G��+��"��RT�Pg�ĂD�� 0U��g��%F�͘�O~�#lٸ���I�8�~��ơ��I0�q'�Az2$i���d�q���)褹��s�̪�{�}s�~��<kΒb	��#O]��&�.Oe���Y
R@�T�lZ�_�Ϝ-:x5*5̸�V�4�$�^�U,�7��J��݄Ly��<C�ct��0B��o�3Μp6ی>���x��o�>���H�)��cu����x�1�(+G,����w����5�����g���#�it��A�џ�D�o�j�Lj���O|�~��-�6�Ψ,��������s�5t�X��6N5�'&sZ(qR)I���P�M���M��Z��'�"����@�[��k���_w-"�v�܎^xA�]:��ayjb��2+�Lh�-�܂q��!��`Ŋxg�.���`dUW\/u�4q�f�j�����7��sgl��Uػw��@�X%]
=y����3� *�m�aD��p�M�L�<�jx�;�3�&d65w,��p�ׇ�N>��G�}Y��Z
ƒ�w�WDhR�H��0펬�H�QE�(uxń�wM�ބ��GJæ�;}q�W��+/g���۷a͚�y���)�p�<97%H���	99A��1c�Hx��9��ˡIkMt�p9�������|yyy�'"X�l�o�F7�h\����q�T�� �(>��B5��4�����A��x�%4�ssKϒ�oo�g�x���S�sǊu�ū�3��Ԉ
M���̴U��N5y���R�3�D�px�z �MJ��_�26���q���!�N��ݻ�v���fɼ�(~�W����<q-I0ԣ������cԨQ����W�a�f�Z�N��;�pW ����lx�/���C����xs��GSk'O+��e�F	�p�D��N`<a2|�[bܓ�zYp�l�O	��WSǓ��斮��-`<�e芝'��?��ʼE������Z��v<�r=�D���N[���ts��آ?��[�b��4@o�G��|E�	=B4���"\q��0�Ha��w�v�KB�%�-�*(,-���@?�<�I��=<��՛o�رc`I
֬{	�w��0ΒL1VFnqR�$���P��2�L��?���b���8����-� 5�P1�k��_6
���;+�قBb�D������Ǿs/��>��Ot.}���ܳ��{\L�3~�3���sV�(���������Ee|��9}�x+�j��٘
�oF�v� �-@2��$\u���/A,m�����ֹKA�� ��J���#�J����AB?�|N�,�Mӧc��q�({~�Kط�����啨��Fdp ��0�;�؍m"�(��ڝ(*�G�/��-~�$�$rN�k,������i�S�qѸ?�i��{�Jl�ib��������-��+��{<���8��gW��Oϟ��]w���W���x�=\E���fdќ�R�Րb�g�T��$R
F��� "�=�y N=gO<[��>ě7����z��_���B�ǻ�:�1�	3�p�e_��Ƒ$��oڌ>:K&����W /��[}]��v�1|�.y1���� ����w`��&8j ��/����zH�"����\��� `��_�bD�?�ԇ'�s�٥>���o��֬�����Q~�Ts��K�������9hPd�����+߄�Tc�؏lk�S&���C��<~�p�	��J�X*��N^3��N�E��:�-G[ڱ����!@�#I^|*y��@~)&$ɝ8!�}L�0EEHdl<r'ڻ!��-��y�H㎘���Q�e�-��ӽ/�6~��z罏�ܗ���ef�1)�S,CsS�]�&=Ĝ`?M>\9W��I�cx�V�ԟ���g��?��{���B��1�\?o�؇g�^V��Q�/q�z�5�=�0\=I�&
�Ɂ'd��ti!iZČw�$��SFz=�OY���$2Z;z��Ð�AL��D����M&���	C�*�� ��^�L�^�  uIDAT>��Ye�oc�;��x2�Pnj��д#���d��M��6Ν|6|d[�q����a*�R�oDc8�HS)�^�t?q�\�p��L�Bbp�~<��P[�G�g�m-=���Ҫ�����ճ�>玅��rV��嫶b��b��?�\6FTI�I��u��G+��[c r��U������,/u�5�t������qÀ�B��`��0�7�`�	>��ilDqq1T�75����Z=�×4jd�Rb�k��&����r��5��q#��.4w� ����cL�ۋ4H�g��	=y�X�K�~͌����iǙue��7�aU��)}2�^����=��_�]՜�ӟ���[f>u^U����p����0�c��\v�&�X��E]*_VË}��$�qѢ�p��A�hif����*T�ֲO���`���	���B&�T���������CM]=�K���Ȍ]�B�=?�7����Ne��-�DG~�p��OG]�(���� �l��(��r�E֫�s�K�5m	>	Q�읱��CV+�m{�{�?��
�?{�6<��~]e�u�]qſUx<�4"�j���kf!��p@� �5����P���v�譔��s �6m���8{�98g�\����8!9���"�1j���ҫ���5�\r	ƌ�Bp�[W���Q,	��٤�����3�$Q���Tח �Ԩ:c����e�Dǆ+�!�_Dӊ �\�-0�$w���6�����7w�}d؁�/����97��|���#u @1Vq'�F�7|W�\��u���(|���ɭ��!��Ǹqg��ɓx��c&�	�P���"�505��,ֺu������.� #G�N�t�/[���O�S	�p�)�V�/���?��5�~%H�α��'���1��q�W4+^!�C������G]�[�����ڿ���|(����?;�_�%��/�{MCI�eye���7�2EQ4K�9Yб%�&�x6�&�7���
rs
���a�	���ۻ�6o���1a�Y8��8�,9ȋ��S��.�5��d&cp���+���'��K.Ec�(�@ze���$IM���H�W�Ds�1��q��ע���TN�8�ٞ�����Gh���(��.;RF�eK�E+Mz�F�2z������ij��|�̏>���3>���~�P@�}~�O$T�qd[-J������d�rlI�=�e�^o�ITN7�.�|f.��e`߮�رu�;�Ǐǹ_,�Ye��a3�B�:�G��!r�q6l؀��f^�W\u%F���(T��C|ށ�h8�r��Lk׮ő#����k�Fe�(�IZ��u����������	(�DB�e[�m�q��X�T��ےi��m*�M�b���jW��������Yvǧ�g�?<���	w~���0�F�?�ߵ�wlg�ʘqc��/^�|\�&JdF
�>���ˤL�������_��e�ې,��
�D�!%]�t��I�����`^v)jG�Q����k�^��7���7�?���Y��o��~X�8n���p��r�����{`��[�v�8��q����m(y�q��Pc[�so���J�(a�ڗq�D4��.8cǎe;R�d�31v#8��i�/M�"�J��G�� <�^z%j+��6��D�<���ol��ށ������I�)�<��w��e?�3P�c�;���6�R,�5q<��w� ,�ՏI����+�u�$��1�7�|���+.Řѣ�LR���8U�<[�@��h<�u�~���~O�~�jT4V�P�����O�Yv����#d����	������2�����ya�>xo�>�ܱ����s�¹��t�J$�&Q)gU����e�A�09�G�����/ĨƑ\��rB��b�8���In��!P$��^y}=�z����W�td%��Ʒu��<�fŽ���&��o}���,�A����م�;�s�7e�dL�:�S�ó��+7H�=��f*8�%$�4֯_�M-�v��RZ�a��������X�� `��߽���(����Z�׏D������u�|�����uW�l��r�/� �㧌���{o�������;�g�N�ȝ:y���ڟ�'2l�Bu:�l��D/��x"�c;t��C�7�4�z�Y��,��q��tlz{������AU���~���h�л����'_y��������?���_��G�
��s�v�ڹ��ϙ8	��Na� e
4�xz��89I�RҀ�믿����u��ѣ�2����)�z��D�<���+/�����TW\}-J�j�tm����#�?�Б���C��M����u���u?���� �n�֭�Q���I�0e�Tq�'�j���� ��.;QHq� ���8~�_I/��"�>v��j�dU9W�=q�_�D���ݝ�C.��
��Z���~���=�����߻b��]��J/�dӑ�m߀w�����O?'��"��k/O��,��e�zަM9Ր���i�0~��npI��!sR;���Y�Q���tu�����MÈ�c�+�㵖����7�?�wQ� �����n�e�Ȑ>-O�v��A���B�yP6�Օ�He�l�N'�f���"�L�%f�����Doo/�����ee\��a�����}��!�U;���ͬ0��c��1oA�z�tN�����>�m��O��5���,���OS���'O���N�A�Ҙ/ͩA��
�S�b�v&�g	���E���2�O���F0�ΐ�r�i�/��B���U�tR�b������Ͼ��}K�_��_3ȟ���f��>c޼�_�Ӊ5UW��z(�J���(Y�v�w�z?QG<�R�G�O���]YÖ,��etH)5��]"쩿�P�վ��N��4��#�۵�Voxs�5����ox��7=�x�	g�:u�iו��Vy-��r��.z�auv�l�!�l�U���h���g>��0*)�D��K�HC+���I�j�͝[7�����ߴ�����߇v�_�I~������^o�#˾"�?�#�!E�Y�H��J�#[��h�#��fڑ,;c*��:��.�V����"����r�$�VlG���H�eiۑ��d�	�J�D���~���ړ�3�V�z��|������������?��C;i�T�    IEND�B`�PK   �X�G���j  sk  /   images/81ad8fcd-15e9-4bfc-86b2-1d5dd79993f5.jpg�zeT�A�� �����e !8��,����<@�������l|���{��ݭ��W�鮧����s���M ���� 			���<� ��_���x��������������� ����1116)�2�7�o��_֣�b��b����y��,�� t$~@>2=�2�s?�  	���Ջ}���10������_� �������B�JH�+�H����_P�ot��5=Ě�0F~3�`LR2r
&f�w�l�B�"�bd?��+(*i}�����70���jemc���������=4,<"2*)�GJjZzF柼��¢��ں��Ʀ��޾�����љٹ��ťe�t{gwo��������5�q{�@F�o�?���y������<H�<��$@A��}M(��f�LD����}��~M���4&	���� ���;@��_�����y� ���^�L  ��D��gV�#���2`E�r
�W�V�Q,眍#����	�0ܿ��'���IS��lg�r���$��5�F�N��.���T+d�U �n}b�B��?�����zs�$�J��P~����$��{$�v8�Z�Ч�:�<�����R���t���=��ʵ����|l�u�,0U�yBI~s%o���4.W3'���a_��l�����&���=E;7sK�V^Z�#�����]$<π_v�� *���cK�{��i��ֵ���n-rx���F�o2�_�x=P����T�����4������b?��kG�u;�Y}Īd�t߈���0��.��31Q�65��@H��� C�Q�*�ݯ�c���M���khۘ�Kig�g�&$��7�D��A�R]GHO?���0���r��;ѧ�����C_�1 L�O[��Mn��R������dD?�� ��d�Do|2�a�̨�<0�1i@͊��>Ccw<'����cª����t��4m�Eu\��^�U�>�"Qr�7Np���I=�p{;!V�jPGx�ޑ	_��P��cq�����y>�����G�O�R����$�π<.�{���3 ���G�R3���L�����l�����~�4�lyv�p��!�����ZF�w���c�=ShU#��+�d��������� s:�4٦�o�dmR�6b��k��q��b�ĬY�栴"?7�">Y?4�W�UzO��#��%r�["����W�eM'��C�9��!�w�F\D�:�v�X�������3��'��b�7}=eZ,IYQ�f��"ķ!�'��|]���mIȫ�+#� �	�Pm<�
���E�����^@I�T�y��Ma�<�;�6>yOƞ�n�����3とߺ��N���N!��o�+ҟ�sH�˺`+���~f�g���g@Dq8������gf񁼓)R�� -Ɉ{�׎�h��z����B�/���M.<�WU�!��xI,�H�6�2i{�����\9��n�9��WJ��b�R*�}5�~��0�T�y�o��g8{z�9���pU%"��4	Pl��p��5N���>G�'I��j�Td���!�@��t�v�M�gF��Dz�"*5�{p7���JK�I2c�_������}Ж��%���]Uz�l ��e��%�$��>�q�n��V��Y��X�[pt����y��ƨ|�'�}��7���ն�w�!i��W￮�vrt�C9ĕ4R�)��0"�[����:L���Z;���'��'J0����1���i-n �K*��x0���Ժ�5�\�B	�t%�U�)�^���т��U�0��.��t1�5�p������F��P�FR��Y�K~�Ms��(D�K�q�V�v�[;1I����ž��F��*i��!�J����.�����X���p��pW��I#�z[	�Z��c�(��`�',C�\�N�����'�����I;�����B~DV��-��5���Oe>
]j��6
%4L����`����F>21~`{Lgש�����9G-��I�l��7�$Y�h1����G���,�>���g?N@[.��h��T�m�D�c��^��@,�JcMЫ�����s5׌;ɫI�y���^���П?�����r����Sq��������/����z�>����(�{/aGI�{x� ���~�%���7�4i�?������UA1J!/s��0y��+Ū�c򗒀��H��E��Nk9'��~E/(�.��s�p�'d�[ D��{��u��jׇ��tL�R>E���(	�2/~�,��r���u+k��	�8�N�}�ǳ�3UD�9I��s�PKs赊�E޽���f��9�F?)����GF�ˠ���O&811�?uq��T�(��{��tT��5�2��I��*E�6mv~$�d�"s�go�iR$Ұ�A��i�e���qh�K�.]Щ���r�x:�O,��P��k�ƚ��߰I:�N�I�I�/HgF�Q@�3*�?�R���Ģ/�G"��ׯ���5�s�/&�JN�t�5'n��͈�����.���(�]�|��%?�i�O��� _=`Uz�����\�w����|�?���ŏ���<Ehn�9w���e	�f�}+����z%���]�옽�����<��fE�o�ݸ�J{jE�m��wpF���"�9�,Z����Y�#tD��Z:�����a̐&?�<зy���z)9�8?���:fn%�0�f��/rp�)
��"�7dP�E�"���@����op����u¡vR�k�VR�4�t�s��-f#�#��Um�!VX��v�=k��k��bJ�J��ș� �ӈ�- �r��wR-�
3J� �W���n���0�Ĳfg�G.&O�p��hT�)�� ,��F�?����Q���
���qw���Aj�_�U��{R�4�U���*b[�֧�ٍ�.��S���yWD �-�m����U�d[\�*s��{5j�?�EE��"z{�?NF���5Ɵ^��D[f?��j�.
͆e:'���C9Y4R/Fɕ���^��=�+]�F^g����yo̰����]Bz0pDuC�¼�M�q�P1�rɖ�W��RǱcΣ��/;M2��[7��O�1�ǝ8����x��bl����ν{������A�1�A����~�1!�Ű���d�s�&�5x�*%�!!��>ԥeЫ�dIh�/G�m�-�Á�ǚ׿��ؔD��f_|[���g��̄�U��U��#�W�#��)�$�S�F�<��
P����\>�
�E�>#��� U���4g����Ls*������&ӽ�8$|�\��;�1��I^��4T��ԇ���䄪�ɼ�rn�B�������*Q�����j�r��c�Dm��h�oc��Q;Mֈ�s9���B�*�� }��7�O1��T4q�ףp�S*�T�e>�M#�>������i{���4u� έ!p�Yv�.��zd�f�}���?�B-��wc������� �{�����qj��P��>�%Ĥ��ZJ��q��;��?�+��I��w�Dc2��YHbN81���V��9�c���79��׃�%�Ux^�z����O��F֭1F\K��h�us�a���e��r_/�t�A���8~��!�A~,�[�����R?k�����K,����юvR���G�5f.��4x6�6��D���`Mx��p\�q��O�6g�)�^3.�����%t{������-kڐ��s���q^�Ώy�����	T�4��\�G�.�kR7H��3�0�"��N/����A/@����ҕJ�ߏ�2�d�� ����������D0�2��/^>Lk�M�Qu䋍�v�gU��f�M�,J���˒o��s�Z��Z�S��y�;d�GYSy��V8TtO��;}���g�]7S�(b1���U��hJW�]B�I���τ� DMƑNr��u!�D�1x�Ys�� 9�8N�eydD�MG����7�-�"�6�+�2�����;�:��_⇐5�W��^����)�3�j:ǁEzy�+s�e��w�Q�����wҥ�?(����ؗ��&UOo�=ⷍ0u�6P��6Lb��Z-P@�	�X�t1y�)m���tzk^�U���h�ҾR�
[�h�ƻw����J�;�}"�]�˅wt�(*�J�qM0}+:>�i���q�Uק�A�N�"�%����œ|0��:%��~�x��NM�4��F��y���_���Tx��u�!.��N�7֕,Q�6��:W�`�]V	��9��(%�~�n�n��@G�*I�k����L~ U^�Uei�(x!X�}����I��#���`����=�ʧ\_��x3����Q_�<�����W��nJƔ��uC���>t�>pڰ�_���G�T	 Im4�-� ��r��QKq�n��E��8{va�@��6��^g<W���'��?|6�7u�iϱ���xF�`Ae�H�>�ʇQ�)/�D�эG�����δ�!�� �j�9�c�/LrMg�5gޘ�ֵE�a��w���n��=.���Nm]�CwߧBz�Z�:�Pn�P��˷_w�\��9cϜ`s���v���ˢz��|<��0v�����ѝu�&8�b��eQ�_m|}��(�g)1\*����@0x>�z=r1����Қt&*+~�d5$��zG_~�N���y?DK��x/�a3����1\ܾ�7=�
 ����~Yl�_H�Y&���+n[��/�҄��c���Et)5+;����u�h�m�0�0�@��M�n����������o�W�Y���!�Bx��_�~��r�?�|_i�`��̈́��H�رݪD�N��hM����>|2y6����O=��6�oh����
��]pe��"�b`~_d��p��lU��͎z��.��V�m xs��z� �aN��R�W骴;��ND��Ն}p3��C���:˜y�޲�������v|����I�Ɲ��j\�<�[�6pG]LӐ��U����1gYb󘦨��\�93Z��h��K�!�>�#�T>f�V�*k�x����|I{�ɏ��l[J>%�u�̚[��4qK�6�[�«��Qo,��K]����;r��X����L>�]��K��{`��p����zό^X�����S�z�]�d��B<{��/��Ӏչx��e��2�լE�D����|��[��ueݖ].v'i��3��T�~]��a4n�~�'���{�7q�E7��y�^�jD��k�-M�yN��-*.�O9���%2&�{&o�F7�9>nf��=�����-=L��Z�h�����M�9hA�l���}@4@�^#�8��W�	&�-.������B�1� >^�>D6�~�K@�nM�l~|�5�a���Va}��\WMbGw�}���K�y�<�����%�A�-�C���ͻ_F�~6�mk�b���X�i��l�3�Y8��#���C�^D �N�L��Lgg;7Y�6)�\�IDo�Ri�#&UVl��Y7*l�B��G�رG�I�F^5=E���n|,��E�k�/��]��T�#���m��{�J ��+1�&ЯE��C�z����J	�<j�WĜ�Z�3#קΑ2ģ�`�lY�7����óab��zF���'�^4wyOTB�(���V�Mjt9!��[�<_�gn�V� ��-긂ʇ�W>���c;��L������'����\�Gq�v$�]�a_%�w©�}�g���	ν|�	��֛��}3�0��O\�;f #�d�-Cfj�-���:�-�%A��9�.��DȏV���h��~��ff�`ޣ�tN��$/���5���B�Oٯ�:I
t?b��?_2�O�^����=�_j�1N�R\��x�p���=�=�DL����7�/��N"U���1����)q{�=a�:c��$����K�I=��?��Z�Y��dK�Ք���Ax�iM��P8���s��9W�4���U���<ը?	�|�K����EQ���C�{�Am��Z��AqQ�z�w�����K԰a����P1|�@�'>���3 d+��O��t���ac��Sŵ��-��EE�2Gê�֙.F6;�����Eލ�_&&�}�K@ubvL���[l	���,�J�@%�px)�֠���y%kιS+M��>42��K�[�18���(B;ں7�8H�x��vR"v����h���l�	e3^�����c�v��9��HCDyO�)�-�t�3��m��(���#嶳jְ�V��p-n#ܸ�t�׎X���Iƫ�l�Fb'H2�=D-ԊU|͏��^ɽ��̜�M�� 0k*�o,�}WzW����������0���e��@C]I\�^��|�#&��O�>��#�KW@��:��n�qo_����5̱&�ܳ¦���s�Z��������s|����GR�������ЪA�k�XF���g$�M�רBz�����č��`L��0�0��hV��U����z��j�0�G~h#����t����O��P�X'�5�j�h�d�y7�ٟv[7FB6���/��]�}N\ߛ�*����izK��u����';������u���
���3�5>����Λ�N/�Y���z%��KѴPx���Ɉ��s�A�
F7c�-�����J	�?��k�m������j,�>����*�@z>�n�yOx=I�Uy?�s==�̝
N���g�/�Q����b���SOUὣ�%��Fx V���1��T~��k�C�b��e���E�;,=��i�g��e��_O�&ܥ�&�ه�bEQ���D�>�з���d�������L�H�@��ڊ�K=�VC3�f�Vf玸���G&��j8�Ά�#Wʨ��7w��.�D������5�V8����*��ak|�x�S�[�{�T���&S�!��/�o��z;g���د�#i)�9���!�ZYR����=��YN0n:���X�˾���QBRԁ*� ��ǜ��Kb�.n�����G�A큹�x(}�*�$��R�n�P�(�̈�p��L!xglC� P����|�����<��vը�L&�.4���5܆��R�뱹xcb�+�����2�ԟ���[��͒g����?Ng7S_�)�F�0�Q��g@�hg�c�H~�G�cV�o"�j�)�U/=T���y�����N����S��*͑�&a��?�M�lJ��ZFE9}v��얫J���Մ�+��䠶��_{1�ŏ|�)m���!+���dW�y���n�U��v��"���eF"ԛ;���0ud�ɏ��姎���mq��>l��J���f����D�{muWw ����~�mQ�>׼�SV�f*)��5�'Q��жWwo������_4i����^O{�0�G* ��K�+b�1�V�`��W]��bh��J||W�cod�)��{���ހ�\��,C`
Ȧ?H���[��͇/����MSς����\E��8�f~<[����ۘǅ�ĄA7����s��JQ����5Pb��Xc-�k�44}�.�u�N�/(Ǆ8��W����'�t��s3�XߑG�4S(���s��s�f�fF�/Ί�o�7M"+賌ak���,��n.�ȱmc��E�l�&�t�����&�yE��[�.U�,5?�q��u��@�%�0�Y���D���Us��p��?�CEE�ڭR�Ȕ����3��Y��^���ɾX�[�@�CG�t
�Q����o+p����z���;�?�����h��P���b�U�u�9dc9�K�DC��>l�<}���2׾k�"K���p�dyc��+�+W�Y�aq�&�ȩ�?䒴=��c;'w,|P{�8׻��-�[��0��� �)��I�c����H��c�1�ڈ]'�z7�.�D<�̕��H��td�A���>���Ui �����,\�p[�EפW��.���}��y#���/!AS�ި�'�v���*��.�R���[�i11���3g�c��f�v�T�����.�|�xj�=�9��T���C��&��XU)5�]�'y�U�qt��흷4
�4��i�j�!w�v����o�7��Y�e�Y���jQ�v��s��b~ �t�ꜽ�qĭ�>�a}���Tօa,žr����ׁ!���g@(��oWxX���?�g�#l�D����*�����h�kzA�x���pU�n�����&��N=M�_Plڷ�Ý��\��=��=\�K��.ڜ�K���>X+�Xz��*܆������5 ݦI�`?:[����J��)ꯊ�@�5� _��D}8�����q���X�����������åq�<�"��.+�R� -5͔ޜl	���!�Sn�:7�~�O|F�4��ŹE ~ �Ӏ�p�����	u�!�`�A�u�������E��;�M�J�g ����Q�:6B��,�����Һ���	/;�]��m��[Es%��A}O� ����]��/�G�՜˚lkIN���#�S*����;��]�_�;��y!��ޖCZ��A���](Q?�,�վ��С���P�YL	r̶�<�5��z�m���;z��:�b��y�IHN(;���&��ק�|&��ۘj�M��`��(��(/It�5F�YmW��>f	�?0a)�ҊRu8�5M�Qq��<.[�����@Z�/�߇�e�rq����R�ɓ���"�%]��MOr��l��Q�1xW)����������9L�_a-9�!��ohHy�=�j�r
��y,P�ʛ�;�^I�)������f�
_u�X_f�U�X{���U8��.qN�~���2�E�{���>l���:�A+���3�Ve�"w���:�͖S��1��(��`���X�L`��tg���4g'6�!����+t�F���m�#��(]��_k�����x�͋Y<��o��9Y�����j׃�k9�W'ʪ���`�<F�����E.���6jl�y����~�{q�3 �nP�[��ѹ���DC������dׂ�6��]��,j�~HXN�%gN��`�Gq2��ꛪ�U�"���$w�?��	7�φ��\��O�ܲH:'���,��T���_Wp��k�1*T�I��o��ف������<�8����d@G⎵�Y���F�"W�j!}i�W}1� \���.��7)��Z��-�:p��!k��tW�)?���㿑�M]�s~8l#��~l*���3�Y"���g:�[��ܵd�?o�m%������]�X Wb���x��g�����f=xrǤ"�R�� �6����<��&��&�����O�1�궓��pL��1,5�L��w�s��+]/;��9�5eJ.d{�x[C���F#�K���s�N��u��W�yzl~�~o7�ʂ�1���x��m��g@Jr� �A/� �l����<(p9�dE�D�7i�cj�*J��q����h��N"�d�$�k��Awu7hef�n}�S��<�϶S��6��O-e�à��-���6ڌOYQs_韦��"�����T1D���z�a���k��?���}���N���f�#i�)|X��V�½P��`9�&�90���+rꢼ�y�yG(X�Kʙp�T�+G�,ǉ_��� ¡� 9{�q����[)�<cV�,��>C�X��ny@7Y~��d���4g�;}��W<g����Vq�����20v3R�"Mǯ�:��&�"C%'��,��y�PO�vǯ�����쎯"��Z�6�ͼ/wBG��tQ�9/ۖk��{P�}@݌�H�Rݒ��3��	�cKh�x� !��]��\����
�];/7�=����'�!?����ͮ/U���h����#�Y?=S��U��p`Q��0�&���Wv`q@�M���̹�\ ���	h�i��Ź�
z�o�mP0���M��MSyl����L�&�u�+�o R,�#^9����������֦v�ɛ�T���G^S���:ye��-�h�F�M���=9�aQ������{7:����|{�ڝjJ<nS����Xgd��|a �+�z`�<����Y�U���X�Ȱ���O��,.��mot��;:�2��@���I?Pe%j���6�Vrn ����5��X�` S+ʅ�3qV���P$�^�<�rD8�-��-O��`��܃����2�W�|S��]?�����R�~h#��L�Nݽ�r=�؇ՏeҜ���Żۻ��}����|���2��7�T�N�(wMN���/�GJ��7ͳ󕧞�ȞK3�#K?�n�4Y%ߏd�Œ�}[��<m�<�;��D�@__��'��e*� �Θ�B
����O�aj�ue]�rg�Y��@�gӬ�Y3M��!R�Su�Ϡ.�x��oh��ܾѼ��i�R��U�R'�)�K�)���un���x�C���A��7%�Ri��;��
�X����GwN�{��L膚0m�7�������j)}��O�Do9�I!�gePg$�;2�E��[�a��K���N-��ʶBa �����+�F������f���{�I��u��o��:-,N9�-u�)<��}�u�d�ˊl��p��^�V~ݽ{Kܣ���|:��h�Vi��BD�2x�K$Ms��ҋ�~o���cW=Ϯf%��yS�Ҧo k��-�0�ڰʿ
YU��͠Od�5cr��9��&�-�-F�!���u�L�jL��]@Lq�V����gރT�e5 o��R�.�Ki8�6ݣvT�ː���)�O0��9��P-'�_�[F=1�H[�� C����s�����:k]�2Ή6��o\k]Q)ﱰ�ˬs��ױ�'��9x���ל��ȻuRG�?1�f��S#��!�3}Z'_����e
nX��'T�7(��`���c�׻ڱ�O%�C�I��������.����E��{�g�Ί_��1$}l�3���=N"�Q&u��Q�\���W��֏NĀ��{_��^.2�w��o��VuaC�B����zբĔ�x�b>�����!G�a��ZBp�Jѭu��$|j�m�nHZK{���{����0�N�ofmE�	�.�r���W�"�x=]�yJ�����r�o;'���4_���A#F?��V���8�hK�\������q��g�F���Gx8��v�=jb��Tdhk ��h��!wyC}�]�<�涮+B.�QLєMx*.Á�!9`��[/����.����$��8:�Y���>Y,hI�21*8�����-��Zݮ���t�����(���Uu��V�:������>��*���JB���^:[�;���σ��`�N*1�ۣ���'���9�_Lwm�g�~j)�<%���7��y ���M��z���$�+߳�	��<��;w[Pu�s/ed6�N1�П2XvKNh>��ix%CS
�ʔ���B�r3�jbg�)B�<k��']c#�Y�úx�x�g��5�J��R�)��m>T��L��#(��ɇA���Y=�sƛ4ҏ(ɶ��f��ڞ\
�]�fu��.[�u�E���n��ukCy�IB�%�fwZ�q�Q���o/��vS�s*�`Z׼(��O��_��x�6^S��LM ��r�:줅�5�0����n��/��0��K찂͛��VA�q����>4��ܲ�h
�i@wZI��!�cTq&�r�ۉu���<��� ޕ\�����,��c���|A�F#���i{����L� ��ӏ��|2Z�����W���CL+B�do�E�Ӝ�e*X�%���(�5�k�Յ<�>�bRv����S�0��WݜH��]y�ۻ�h=ǥ�ŀ}�����jLGL<�j�0�#s����$i}�)n��.S�oѓ@�1����-��P�>�
��Ϯ�=��\c2��_1*g�f�n��A)q�9�p#���'9l/�osr�fs�.�[�lO�����RY�dH9�Fb���l=ؼ�A��1��m��9�k,2��d��l|3}�O �βɜ��
��ӭ_E]��Jq��s��H}>Ez:�;��qV&��@~;�#s�p��*7�L���е0����%rͫ[���sŠ����R�bj�m|�]�FwTb�["U"��0+�@��h�gܽI��=��x �D�����d�QEeћ(���9F��w��k����BD�(���K"�4���QI�.�I{2�S�n�V�1/Ã��U�߃�g�UQ�3L��/�������_�b���`a�W�s�d649���?k��'6ee����w�q�*䱣\uy
�?���G��EN
�R��s|}��'9慬9�RiaRo�ů�6_��� �2ˬX�+gX�a��X(����m�T(�;���V�L*[ ��� �H�7Y�5dݤ�h�c�)�D�[�9�a����M����$��H�@ �d�^�8Oʿ���h5�}4��gSv����W`?w���M�-���	�q�i�HѪ��޻�X�tb>LfG����^�
�[�����g ,3b}[��=A�:$��4�zJ�� ��)o]�l(/,/.�^�D�px���/*��-T��37i\���ի�.M~�K�����ÝN��N���[2��*fl�?�� ��jܣ�r�c����F1��ߍָi!�L��Rg�2��Vx%���.E����������4��fH��|e��~�^HV�!�c<��k�c醗Ԛ�!L�ڶ��&eW=�3���拮,��_�-��VP�B�v�:e��pF-��ۭ^IWߐKkӈY��^#OwA 	:�5��0��ub����\�қ�7�#�N�6�<\��px<�u��?:>�� �Hh���ٯ>� 6vJ
�҅ђB�����vZ��Dg����|�J_�!����=�����xE�����&� �on�7^�+fFE��l!�!����v���Y��2��3�U��r��:|�,EF�ۊ���o���xo������f[uc�@�!�������JM�':6�y��ZW�3˞��ZG(�M.Q�0�ڔ%�}Zc�2m�$����zgb��������sd�b�qt)b�/�t n_��֩E!`�R��
�Sث�^O"s\�W)�\c*�w7ͣNz��!�r��C\�Q�ZN����Ǹ�0������5��m��zo���^��
kZ�`��+y��xRx{�Pv}粘� ����<�ξsJQzq�w��Z�B�t;3����G��>����D��]渤$��}
����T}T?���\\@�#��`a�sº�M9����������n�uşqD�;�/�|��`��@n�5�|����#�NPd݉�(��l��ɠ��]��2y<!0)�&@��11���I�@=J�.z0���93'��#���3�n��)nzF�vQ�aGծ��V�G��h	K�R��s�	�Qr�U�Z�;�~!��)���M�%�'n!ϻ�ZCv�S,F^E0��6I�����EHa7f�9T����R�w̔�Ә�����ď4{6���I
�=o'#v�G4�q7�~��y�3��q�PƯ���F�u-�I����\�9��I�pr��%v{��+
#��r�	@Sp��a������mpY�#��Ej��	7p�nB�����w�:-��j���PU%N����zP���C��O�Aπ�F+����P�/#���\���!u�����89� ��!E`L�
x[�������'+]Los�#
�E����N���j���8,��/(;�`�W��"�� i˵�^��3����jj�k��6E���&���1�i���H�6��v����-4
�FC5f�̕�U�Su=s����z�>���{<�x�emq���\���pժ���9�/�L6�)�ۀ����� ���M��:��-��r'��;���O�5�3����π��5	^�˫��i�5C	0���5g+�V?�}��[iD4ަ����
�+n؄��4V��2LP7P�{m����~M���a���:/���0,�S��ܡ���\����k���*�V�4K��u��Z6��M��7w�]�@�I[�{s�kac�TY�$Rº7{�=
*���Ha�qŬ^EWf(�������]*�Q����2~X˞�s�߭\��Cl�"=�����G?bJҞ���p��
�ˡ�i�,Y]���E�X�]��	�پ�:Y���9m��2ȷ�*�1LO�(��C/�[�V���?L��ȋ�K��:���.��0��0kB9��~x����Ի�wCt�񧭽���?Q?�@oX[���CSN݆`�&����e�K}�nsz��m��'�;C-��G���1��%�f�4~���!b��M���~)���E`�*��7K�{��p����3�k.~��R�NV�d�!���v�&��ҡ>m/�`�i,��aד��4��ȳ!���p��2Q�O�Qc��j�ŒdS�;�q�&�ӣJ)�	�a���'V���;��4�k�l�d~��g�V2��
���Ԛ����dȐ�%q���wV����W���C{�:��Fo�C?�VN���QLҫg���Y��$Mݸ~���x��[k�jBi��pR���s��oO��52w2���o�}��迪&f�p<���#5(��%zl�m�Y��p�io]�F��1�R��=�OJ�<?횒F3	������E][���ʊ*SG�/T�JQ�Y�^�����0�H��jXR�iڱ�z).�D�⺲�ri���z����_aICE	� ���t��!4'��<�~A'i�,7�`���;1��Q ��h��F��de�kO��7�3,��&u�����3�j}���C���Jy4��m��B���G��xS]��US�|�g��6�������3 �^��3 Pj���D�u��$CO�?/�2$Iޝ�����U��^��h.���`�u�ORy\�E�Nn���T�s��7x��W�b>�"|��
yʒ��� ��P���əiK5L�[�A�&,���5�}�P 9�~CM�A� o�nZ�N<�Ӥǟ�*�g@��pp��6����n@J;7R��C�@ԡ5�GF<���򮆕g�TJ׮Qi���Ut�~nc��q`�QGE���iA�>��9w�R&ו;�绥אoo7瀵x��B����2�5:6�Vu�^��~�
~�����`;u�X�j~ϻ����s��uu'm�0�y��UO4����oO�P��\8� �>Y�s��/�X��-���e�+'���W�\�@���Lo��Q9�h�o\�ņ�m�ݵ���,?z��j�Wc��o�;Z�wjg��H��Wi�N��ƽ$J2L��佲�%�.x��qu�3�S"+�ӛ������,mkrjN�w�<���w/��l��U�>�.��3>٪4��6���1R*׹���u�c��4�q���*���Yk(Z�}Ɋ�_'d��7c��?�'#����U��pEz���g�q�?{�5T��p'jQץA���Z�˼�x�ײH?y��>e4�7�u����S˹�S��U�@�0r'ḃ|ػ�%�OU53r���e!�BO�h��i�� �)��W^��ᓺ镖ޓ�����t)VږT�F2�W���	dENSꨞuؙ� $wu�>*�3��e$����xjJ4��z�±ڎ�q^'�3h���N���sڞ^����y��6J��I�;����Ұ��Ξ��I�"�$�b��#��>ż#���h^,:q�� �8��/�Ǝ���ھ�3�Xm�]0?.B���
�#��j���_z��~a�vt����J�S�/��7�
���k�8]8��=S���E?��2ɥYE���Ǵ�s�����O��e&�D���u��Cg��O�YkyC#�
�`�/3��R�kW��h�3�g<����!����f_NyϹͯŻ"���b�q�S�Z\�;R��=>�/�����#��r.���~3�k	vc��K@P��j7.�5=�SS{���ŝ������|g��2�3�Ir�9�	���v��{��n�K��*���Z�������u	&L�y��ʥלYY	���T���wB���b�&RL��M_I�����e�����f�>N*�������G�ljo�sd�M�q/U	��#�<�W�m^����x� �M���}�7�;@K�M�➭�w�ߪ����f���lO�'�5�Ig`���(�<,fX�I4J�"O�����~+�ځ'i�	DGǳz?q�#O|����P;a��xv}������kʡ��̰��	��͵�W�vw�����obO���>?Kd�0V�i�r�g��n���d�Xؙ���u���h�1�(��0�C@Đx]��i,QM��]8�Ѿ���';c%䛮iF��]��ޚ·�tl��9�`5̢Y��{���q3���GϨ�2Px�����e�Nji�FW���|�����1���5�"P��j�<��p�6�B��N�w�N�!�#B��n�%��(�c��$J�n���.:���{Y,���<��̜�9s��z3Cn�w��JP��5[
ʍ^������)�`��bK,]E��0v��E+yݛGҨ��"$#^	ؠ����Ѝ<�6�o�4��c��6|�ˢ�IQM��!��e��1�$�+�鮿�/�N���9m���Sl�@U_�[^�����>�to�s����R�s0���l�?͇e?.���_����Ȩ���9�@,1$=X9�Ki�N�c���`��_�$�V�T�uۻ���Ǐd��E�Б�ir��1
��E�����J��ao�FG�����'���W��b���ב�ݼ����,T�G���T��}�|���{��Kz��q�����J2�ktv��B�F��Ďq�[ǯ��@ �.R�	L�Zl�F�d��¾1���x���<'�b�Q\�<���ĢRX��
�YĔ�UBcQ����N�,�c�c��e��:�v�f^��y7�2BX�2GC���9��/�G`�.���4_}��)������K�/�3�tg��rS�|8ֆ� �#ઓ�֨{fL�[cps�� ����S�� ���M�
��/≛�Ӊ�����֭��$� �r������_4���)�,�?�˵8�ۜs�/:�0���Q�h�!Q�IªJ�������X���$�x{��,:a�e�����Ng+b���-�O�j��gʾ*��o�Z�˄��^�祩�e�Nc�݆���v���R#$�߿��j+�x"i��١���~����T��e��R���G�onѹ:&Oj�W_F�`ĺ/K~��T��:�X)�R@OK�D���J�41���|��ptRb�H2�$��Vz�QM���8��E*W]앎�&�FAZ�JCL�\�I����^�z���a2�7��Ǩ���ϛ%N�			Hv
>W�d�L�=��� Շ��z�~L�i�-i����O����5��B���`�w��(i�d�p-�;�U��"5�`�(�"9��(qf�8,����Jf"z�*�O�U�����OI��ڈ���7N
�-!T?���F˄Q���^v�U�#��h�Zdʛ>)�E^�|#�bj�G�9c-�G����W*��� ���v8�3�|��.�����D�� �X���>s@y�~T��.�$�)��a��B���L��1�:� qfi��wMܕ��w��[��Ӂ��%P��u��%���]�)�`����ĉ%��7N��XC�vOM���)(���n�1�����_��07��h��z�z��v�(����gQO
Y����[NrXΩ=iw{?u	O9`������hb\��Yڤ��0�JoItT��U�xsڠ��"X�;����U��ޤb�61xRX�k��
ZM,�*����EHo^'j�L����u���f��-�c���.8Fq��J���|��dQ�>�Xsf-�w�v�����e$h�����_a*F��w��F!�� oH�}�C[O���H�l�~�gO�N�{�}�Տ���d�;�m��׫�2��g��Y�oV�c�K@�f@�)�����t�L�9>���V�?I=N.r-yS�3���Ǚ���S��I]�����~\���h� ��ڞÖV�1Lu��JM���Y_��lC�a�:l�0�G@���6`W�էp�F�T�����3X�mzl�D�ߧ����\�����Ɏ&=�����\|\�{s��-Y�9�T�6'�q��0Ԇb���k�՜lG��#ښD��ߋ���ٽrt8����9�|�,���!*��9P#�/�ǆ�p��\�J�U/�����'�.׮�;�6��G�W���)���}kK�]�Sl���hc���m[�GEFl_����3�~I�)��ݠ��丸&=&MJ����evw��.?��
��$�
�V5o|~��3^rL�26]�3<�~܃�ש���y=!#M%���H'�>d�!���fa�� �i�
V��\��	'�Ӆ��_�	�1�DXZ��m�m�dƔ-�/�A��|ny��9n�eh��D����"��w,'�oWf�p7�޷V2��-�p��咚W�ЋPv"I� cg�zf)#`E0d԰��?����6'M�Y�#�
��22Yn��Ss�A��f�KW8~�hz �Е�)'�M������=N������Uw��9���`Z�����U���2�%���f�n��_���� O�*�U�l|��U't�p2�h��xW���n���n=ɜ���[�q�Wy �yq�w4�O�����-jQ���z�+�k��kCv_��e��a�w�QZ�B3%�V��&Ħ��cPu����׺��#�N~ \�{ 0���%E]�k����hc��T	3��A�?�$�#��d���� e0���5���=^��=��{��n�ᘫ�,�k���ث!�~�����Er?�%zL}m?����?�/9��L��9�
�X��#�����P9������u�fx��ht,�J��S�kg'K�u(Ԩ�X�cD���r1�E��Sg��갆b����9e�]�w���Ʉ�4���ϯw��k.ou[$W]0,���! xʳǋ5�)��_�롩
��#7LR���Wg�3=<�Ή�Amxv��e��sq����F�k)�bg�a��Op�hl;��j��ܝ(��v�~�c"QVg~/������Kp��KON�S�.���<�FTerI�kZ?�m4+��G��njd������",�����Y��"�a���q�r�l���,�N�k��h�1��Cg՘TgP�����y��b߷��Gka�
� �n���;�59=��W^��IYRߓ9��_��V�=Ȟi-|���\��ơj�W䊷%�64`����>��d$��|fl6���.�>V����EuccF�j�}�)ODv�Dp��x��t�+�Q(��k��zB�'��6KB�Y���H,J$��b��$vD��� 8SʝG��"�g�����4�F��zz��E�+1_��;40��ӓ��ar�z.�A�*.D�
��%�;W��vqC60�[�����'�j��	<[1�@�^��0k��x~���T�r�P�9�unSMАI�����^�zŚR��,��b���i�y�K}T��BF��fL�����x:lXL:�]'ޡO&˳�ƶ(���,S�Q��;(��7)�*���I-o����Q ��=�X�!��c�<��/Gͤsy�z�_���ŞQ�ؒ��8Og��&&�D��J��X��I���I=�ɐ�Maa�̙d�w	Z/�U8	��6:s`~֎���7h�.�����Q5re�o}\������ɭV��#�g˄/T��w��R\ˆ���|2����ɮ�ldvl}E�6�����ӯ��}����˛&sA�f*�g���u��i<�����.ɚ^W����&�D�F���1P�NXrnm��P��� 	�_W	ŗa��K���É��^Z��<��8��2Վ�Tc�]d�OvI��B̤Vi�f��R�W��(�j��6G��mmb�D����xok�
��O=��v�kYTw�zyS�-#3�`u@S����z�����|�V
~a+��h[�2�9����o}�˅9�8�I��K �W3����r�ް�ʩ��WKx5�8�WS�x�O�D�䛂�n�7K6�ZL5;�l?�����-���n�/XiaTjSG
Iҙ���W��r��x�a�zT=Qu
���C|�����m�4eU�&�FҜ��E�L���K�M��K�Y][���S��S�j+�	�7�� ��/�V�M+h� ��d�1u�g4^��j�E-�hڕ�@���s��L��<�������
���Xk�!���r\kFS��OգML�\�䊋�^�P{)��橋�ҽ��GP�ۏ'O�U��h%S�4�*4���|����H�.�1	mHR��Bfy,'1ȏ��}d�#C�?-r̼���<Q��ѐ=ȩ���,%��0m-���kY����GY����)볝	���5��ӘkNCٿЮC�zq�����Xy���i��!Ɍ��p�ӊ�_�|��F�S*��~�3��xwA�O�j��'��5,v.X0Cw ���p7>���t��!�xQd�*�����ya��q�����q��Ϻ�eQbv�]�_���G ��9e;v3�b�\ְbWf�o���]}ROW���}7����K�@~���a`�l�?�׸�"?#�J�՝����� 	�9�� �T��2�����+G=��Q�$���yY�W��n�?(x��_��/�
s��;����:���L�����w#���^���n�G����C�Ӗ�]|�ؔ�Mu�.� ��}#/ܣ[�^~�x|���>:p����R^�����c����?ϣe6-p�E����_˯~��>�����\�R���_�N�ћI�ղ�qF�xq9	�WQA=[F�[�$��y*У���[$J@%x��n�R�`'+�w{W��/��ҌG�Z��c�9�\1�=�\��kd2Z=pp�Ǝ{ ����}Ɵ�P�7�!�d�A���c%b�&6��Ǥ?<[i{(�*�֬?�`�oe�vKG��g��^�CV��M�EyD RN�p�%��j��S��1���;�Dp�>յ?~���||q�	�.S�9=R�����/HR���/�̆.�0V`�A��1��#q�m�N,?�ጉ�b(�d�u�����WB�r���6�c⦹QG�xA����d{�x]�y3̮1)���%�5�s3$:3�L&'��U`�X=M)?,����/�l��߿r���}���2|{T�Q^~?Ǥ�%^-1N��ܲRN`wP�Xgm��o6�S`�� �a'���}~6��u��5p�F@\���Y]ܒ���3;ў��e�x���4Wo@C���Yg�ct�V$3��k�Ϫf<��-��*�S������FƭV�kݚ��F7�Ci�����P#ul�_��~m���o���ƅ��V���?�h�O|��y7���G�͑��£<�=DA�9�|>3B����cZ"��6��!�&�������@�U��ƨ�N��n�ًO���Kf���a�� 9�laأ'�=�P�$����$^Sb��Y�
��yO<׹�/�|y�5/�?do�;ȶ֝�X���w���v�����sN�;�j��^���\:�5��8�pk�S�O�V+0���B�|�E�֣4������Թ�ؐK�`o��k��bO�.ZR�:��G�!z���)�)��Huޣ �M���81-t��x�H��dK�������m�:�쏠�zY��?Cn����Gz���#��{��͂������O��˒��߅R��J~t�Q*��O���qx�����v��Mj�`N�H'�O��3��u1��&0�������e���(j]D���+��-��V���ƈsF�ס�0L�9���N�!���w���挾��ͼ������LE�-ƏIߌsZ��P��Ϥ�0�����gp����-�Z����Kִ`�!�Y�%�_? �HQgO�oA��DW4b#����3j�D�-"�bV���>@���@�$OJ��"n�ucJ�ފd��V*�=��%\ie7����)��1؎OM��II�vM���ݮw���^��֢1L�Hh�s�v���C_�p�K�f�O���y<O���t�z P�1k�9��T=���9�r��,�~.�O�*������1�i�*���[�Jb��2�MK�W��;���O.~i�e�^�ϭ�&��RA:��e�؇�Wr��s�����
�^�^xF����
��k����]��q�w��K���HΕJ���#)+�"����V?�O�>O�+����M�����JRI��H?��']1��=���҆�"��#�7e� �7i�Nv�o֨F�����j�$m���՘����a7U�JP�A�o���/ߒ�΃b\�>e ��h�|���x��z�C��
'���J4	���s�,�]l���j�MOIe͋��L�c\r��9�>[��\��e��ig����5�Zu��}�Ԣ�*2�w듫���AF�l��Į�L0O8�R?��/���|��b
6p����UQd7:��� �c�Ą�j��1HF��\�e'�v�YY��l}ʍ�I�nMJ^��d�YN���o3e ����m���&AeX#�S��)��<��9G<oh��B��ߐ��a
� �?꽒Y��ҩT��I�	�	�o�O�s�J;'��G�pw��V��,'d�E˲�������x��������/y�g�-�M6cV]�B'�c
�u����)��_�iv����7E~)�5��6b�յ!��������3����3_]���b��6��6|��]��.U#�el����L_�:+�o���x���S�8�cԙ09xg��$��.�g#
�K0˦�-vX�O�j���C#�r��U";)������tk|f�簡/=O�0G�b��Xj���x���7R�όL��� ��+YuLݍ~=�,b=á���Ʀ��4�`�.1��;y��O����P��
��S���!�F�NzaF�A���P����zjp5��㊸ �Q:p
���%>g�4*�:�9ї�H�-Y�I�߰K�� �G����>��.��<6�iB��}�l���c"��2?!I��թ����հ�@츚H_� G�Dz�G�^���`�:�@M�ЊG��qӽ�o@X&4��x��:>D��Bޫ���)��B0qN�z
ų��_��T|�a�;���UXWI�e�{D���Vlw}��#��6m��
p8,�9U�� �4�S�0�V��%H1e��C�k#*p��Q`���r1	N����b%7�ؑ�kN������r�q���Ay�-�E��q�_B�mmu��4���b-1��7��h^�I!ݖ��c�H����Fhk�ڟ$�
����֎@&Y�"����&���j��ɧ��lO��-R�� A_�_��wG .��J�8��Z��H�>�(3�j�:$sC#�Ɯ\)�>��P�w=y��y� ��#C[�!��;?_���[R9��E�\q�rh��S�&`����e�7��ӆiq<��!Ǐj�k��}�qb������jZfl�X�1�DyZ%�����ͭv^8�ڴo,> %m¡H��{f�=Z�X�QQ�¾�
[�`�Ñ�V�����]�p5���>�ߟX�S�\�cf�%\�S��Q�}�Z��B#�{#b��j(uI
��2:�ױl�c��$p�^e�	�� �o?b��7�7�j�i�3�jޕ��	��{�ʧ�1&g�aǰ�B �7��\H�i
��,$e���g=IX��8��.ߍ�,� ��ԀtZ;��;��E;���W����m�3�����1�*��'U�9�涙d5��[wX�L�Ǎ���ļ�����GuR��d�}t�e:�a� s��^�� �*2�9�τ�v�vEJ�]�h�|��Og����[�%h0�}��'��5��6�1+����Τ�o�P��~����@���b�4[�~wft6��Er���ά����Cx������յeh 9�lV����{�^��6z{Z���d���7U�ɡ5nh�"�7ae���e�,����̸�A��������1��h�gZ�p����F���x�:b./�U��a�ϵ\�U�:�ƣǿ���?�x��u>�&9�:.�e��H���!����Tw>�"��ՕV������s�[��OvW��=v�e��>��Z��M�揣�t�a?(w2!{��և���u��Ö�]7=5�x��k6a���ߣ�U픺�B��?�� �47���	���{�1�|�pO�4G�ڦD̏WY�����������P����4��������c����de��<ѯ��Z��� ���O�����t��V"�e�b�W�z�C���"�\Ϸ`�E�����j�Y�K*[+�T�C��{���v�@f��V�Ha��4�U�"�������Z���(�����.���W%2�~����$X ��y�G�ǜ ��I�W�}� ��[��Ύ�Y݋�-S�0�2������xE�#��+��y��ٙѱD�c8�h�������@=��_��Y+�-)����磱�'�w*'��6N=FaF��E������z`3�-F�s��a]��T�א�U5�Y�����%؛):�0a�E���W"��^Y}'[HY������@�Q	J'�(�4��<�x��_S7�*JQ<f��-!FL(<������{���{�jEn��nj�/�ɞq��5;��'��`ק����[�9�X����AT���9+��R �ɫ�71��߃7��Ͳ�j���
J��z0�~���v��ӕ���F�9����Ŏ�s��5r�Ad��\<�0Kod(.Lf�C�B4P�&���T���`ր����`�ӯ�u	�0u%�N9"�9~|�CCC�{[�������	�-�����O�hh\�7�cZ*��f|�ǳ���_�~��&1��a��+@cx�`-FV[T}�=R֯Ym�et?s<�m7k�7ב�댙������������'/��L�d��K���������4X��zB�����;�6��uD��^>��H�b�d�S?�L�̠,@�j��g�.!po�U��|�a��=��"!�~Av�����& �x����,��>.O_%D��j�ۄ3���~�|��"S�*�'�:^E�> Xh��D�Մ�^1�]<����r`�����F(r8�,α ��#G_}�ֻ��d�*dz��Ao/5�����0H�Dx�6�D�J/��~,h�7`�\�4ߧ"-�˦&�C{c����X��R��BY�m媱O
�.��{&�������iD��޶�����t
@�WYR����Z3�ۉ'xgV�Yߒ����fh����Wsi�&l�f�?u����#��[����ɉ��H���D���w�f�����\⊕�M����%�};���-�;+)�������}��t�V�2��Q�|��7T�EI���<�q2�*�qכ�YS�ˎ��c��g����z58�AC��T�/���X>��s�E������0�EA:vπ�3jB�[��٨%$#��
�W��� ^�9�#�X��%(�>^{�W`Z��,�,V��"]���{�2��
�xo�['L7�@p�.�S7��#X4~$�ٵ�0�u�_I�ͳ��D�*�XIwt6����B��Wu�!dSǐ�s���6X���2���9��yYQ�s�������Б0�_Tjg�4�u���1� ���d�FޥŲ΍Gs\�#�W_}̘��h~��{� ����5g�H�\���R���A����HQ��\��'Y)���p��큕�+=��/HP��< ���#	�p羕K[��0�S�6��S;*9]D>�|��2�|��u�Ix?Q��į���-�=�cs\��?#8��Ccb�n}��]�ۖk��m���T%���$�"�WP*�c� o�����(p�X�s� �����]���Pǻ����NIo��Rv?�"[��_{�&٢j3����ZԲB`= �K�D��֍��ff�5�_� S�R?%��PQZN&����&H��+5�����;ۼ�՗�;.�Ec~�N���隑�Z���F�,1�]DR���7ˇ��hCX�(��[Hb�z�V�C��Z��iA�ldcjq4�(����Mi+Jg�_����b�̮�F,���%���#���$'��"&��	Y��73�	�uF�IN���뭳L�������îY����O��},���A�v�9h6� [� h#���Ė�n�\KR��X�,�r�7�(���i�8�J�
L�"�H X^ay<�f�h��ag9�^�P�qvW�f��寉a���e�T�^�)���
T[�a�W����P�tl���Px���C���M��G1pw�,;QnCx����N����ЙS�s�"��.�A����W��dɟ��������c��k����%��\Y��'����X�J���h8�s�oH���R-5�%� �(�nߌj*�= b�� �s�h|Bt�� {>�^�D�<�rq�'vq�T��5׍����Q��:�> �ʽ既�%XX���`A'�cj�R��d� |�=���`-i��w,����ς�u�W�d~�#���=�_q�v��cM���>e�y ĸ3����^w�#�^�c�
r5}���؁��;�;�zRn��4l߰%�Y竌�?EG��0ݠ��Mc~��Ⱥ��v��1�ȇ��
u?s��=ɶ{���j"V閑�wN����k��p�jp�g��h�[����kX��8�7��#���B��#��(Wn/d� ���pBhI��n1��͜��cȕ�R~�=����ϖY>�4��k1*��{ ��8m�Ԛ+����> (?,ѠU�L<�y��L_�O]�{ D�~`�!$�����t�'�w�$#�_o�֮@ ��jv%�P�8��x����5��r��gOY�b�o A� '_y������h��y_��1����_�� �cĂŌ}��������<��L��Jbf��W�G�wA�]1���Mb���.:��!#�0��_��{�V�=���>��/�h����<�z ��wx!.Z�A�� (n���N���*i��߷�<��PK   ���Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   ���X?S��� 2� /   images/99226213-8268-43da-ade8-d9d07cfcec9f.png�gP�Y�6�3�3
(���J�80�d$g��AR��!I�,y�$9i����LJ݄&������y���s��rW98���k�u�k]k�C���.�\B d2O�VA H���$��̓�_~u��Q#�7��+��w|��@�� ���f��
|󆋔�������DrX��8�<w4�pp�Hŉ� �2��架������ge8p����9~�����9~�����9~�����9����D�a �6a����s�?���s�?���s�?���s��W��
?���|���t�+�p�����q��ds���,�r3�A���7��vaj�(��%'�	�ψk���XRKj�^ی�����~��Gz�޼nq�"�s�lz�c��*'��B���G��*����'�t�����Ð����9~�����9~���Fy\G!�~���AN{�8�֤�M�,�-�U���0/��w�Dd�-�h/j�`��z���L��qe%eP�Td6�`�$!{+m��+�H�0/0�EV\&.1����2wV�6Rer��t��=	���n8X|��^�V����ϕ���-¯%> 6#�
{q�$-��6ﺴGDW`�3�O�5wr�~�;�VNYv���.�7N''kg���}��:�w4&vy
|�4;�k��:�[�$���L�Su��u�w�4���Yz�+�,$d1<�nە��f�=*�����o-;+�s߾k9�����#����0I3��\�#n�-�1�i2E�=�]KeS�g�~Q���z?K\���N}��N.'�M��x)~M�銶w�����2�-#�z!C�܁�����k�U�<K���5,Oz-�e"l�k�xͦ�ٻ��Ǐ�U2�+u�D��uLǭ?U����{3Go}�5$H��67�Ck�g0܆�����<�s���?H�&�����i��rJ=��k���p��ҁ�Ɇ߿Q!aYP+ڭ�ұc�����X�."ί�b��$��f�@�ى�a>�[O��w ��[� _7+�����~g�EG�+�}X��$�qf��q�VB�<��C�����B�o����Y�xj������g�bh����>�ޓ�̧NLPK���ߨq�nd�����B�[F,���O����o��)<�j3����J�-�}^3�S����q�o�'<}'�0M�F��`7�bqmwi���~3��քQ���dFK[XQ�����5����b&��-wd����^H8c�V�g=m$�,�l~��"\D������ӕ-��/Cny6�*�)�O�|�����8�??~ZK��ɳ����[rm�2�#i_j>���1wY��l�[8W.5���P��D#熆�L<������"����Q]��]s��蕄\�y"���;�˰��G�v$��T��Zۭ*H_ݥ��<�>�e�g���P~8FoY"4���i�ɚ
�29�
��g�'٘,�����%|�}��ݙ�F�k&�{ټ
/���\�.���� B�v�ώwt�m.���v���2Ln�E;�3&�e��Y�zDU0�GѷX��R�޺f�&�]0x�;S��>	,	M;R�v�-�)�Z?3����Q��Hs��H����
�y�٩3摝je��4���%{c��E�[::4j���T�/��~)0���o lC�{�݌$O�4{!0uUe���1c6�s��a]�Z�~{0�X�����,��M�4-�F���z����;�N<"O�?�4�q��|�ɗ��Z�+у���[��*�������^�Q7�~����w�㔭�S'����:�X�,�����������K�b/~0
آ����nXn��z><Sj*<�Ij���}{��J��⃖��.���C�\�r�J�l��2�|�-5��u�I�>6k:��y`޸?-3��׺8;K�{�H��d���A���G˝�����ȩ>�ZhO4�h!5n]b�ݫ���R�4�W<+�Ej��7i��BS9n��;xZ%�	?�8 s�<n�%̝oz���(��-��J��/��jX7Z�����(i �_N��Z�û����y�soձ1w�7������2UOZH�N�-�Z�G�(6���oEuE'�pu0�*�S?�=_B����"�/FW=����ټ�*x'D}�}�6�
�����u�:�j��:�lГH7���3Hk��?V{�X�pEn9p�-g1���a �������5��!S'�[ԗ��<`uy��mZ����ݣ�<n�LKǳb��c��`Y�4=�t��?�����>n�~=�-?�1	�/s`|��R���x�g��i[k�����h����__�J�U:ڀ�z�L܃��._{�(�%'^�� �N�c�e�ڔ>���©��3p�B;�,����L�:6h�z���"�Qy�*��hu7r+�Z���y�6��s���Rv����Մ��eܹn���Y�ۏ&�>��[M�L�T	8��J��q>�x�%�ɦ�lx;��ƙY� �ZR�pf�u=wR>�:	��l\�����������(����`!�x����s�Z5� _*�ȩ��@�a�=v�0]��0�-�7�;��ձ�i�&�6_���<�Ik+����>fͨ��ѵ�N0CBK��R��J���j�u�X�N����{���R�6��t����`�g	nK�3rT]ݝ��B��6�|1��`Ba����9Ob9o4Bz�5b�V>3�s� �8	�c{7?�� ύ�b��.�l�*_����N�6�~?y���nTy�/~�8,'i<#��Q�n)��������h��ܖ���7��}��c�:z{��$6N�����:���g7ŎU4���4�}	M�M��f�5�����S��+��pz�e�� 9��BEؑ��#�*@hL�N��o���M'���E�e��h��$����0!���d����}) n�+�~�D�is�=`x�� ���q��$ bƱb��4���/9�0��������`6�������e-w��俀��� Ä1Koc�r�o�v�T"5>������?v� @(zP,{��9�/Yw9f�k�:ͭ�V��H�}��9�Y�o9Z�t��=� ��q ���[}�0
)���|���� X�E�������ѵ������M���Av, +J�X�<>��zFk`jF!(o�ӻ�U_;�����6}�`�p�=�5��e��������؊w���ǡ�����&����'W�Yɚ�HI�:r�������������Իk�oR�k�[	lJXN(a݃���-�������_<V��(��Ow�f�b��g~���ٗ�޷o�h��j�����铆�R�+k���)E��0�GwU׫��<�ݹ���Yh���.Gu>gx��l/���u��j�$y��h�����S�gE D������i@�V,�(��8,=be)���]i_Q�˸��|�FO�������1��U\�>ơ6t,��<;]�i���C�&?z~>%f����V�_���x�f+�,�`�����A`%���Iك~�llZ(/4��\g*�}�~�a]#�1�IK�
�o�z��bAz����P���}ε��1IŠEUUt��1:���0�{Ӿb�=�N��@��[������^4�7r�?H8qpߺ�yZ������s����~�y.�~�y�h� ���!~�2���0�����a&P�so�!l�;qp5	�RPW�hN�>���Bad4ڴ�h4�%ho��r�Ǔ~�}��ܼA������~NGǉi�_x��	C�����  �n"���P��;�Y�th�ԉ����M�!s��y[�y� ��2ǬK���CKF�4�f���ɾ
/��Ryp�`���t���!3��z�{F�Q\�[o�h�(�A��&@�h�*��E����U\��Hvѫ��Qx��0W���z��7!��$t��2���,�mO�����xj�ǋ���p��q=��_��7j�
���S� b��o����@�[�_j��(o8Z�W1 ?"�4#��ɉ	�)�Y��E��<��f>͝�M(-���}����E]u����&�j>��b�}�h�`�r��*� ���~�
dG[���s����'{k�����hvPO��L��_����/z��O�	��wK�D0�P\R����=S*���Mx�vh1C�cܑ��U������z �
 ���Wx����ܽ��aGn�s
��P� �����@���Z1��{x���+.~0>�[ ���큖Ԝ�jWGwynˏYC���ì+��֎������<����jEmX^�J�����d!�kEE-��������A~QD8F���İw�&~�p.��B�� jͬx��� q��E2�@S���Z� q�1sv�t���+,m�@���l~�5{�R|��� U@|��40?��m������F�O��f���:���pi��+0G����$`�ׂ��g���Ϋ���>R�Y�U_���om�MT�xy���]��;=;+�� %Y0fqiCܱ�>A����V�<��P��3�7�mf��w����pg��j�@�i���a��R|�R�0����hh�2�����_w��f����������Oq
A�j�a{l��������}PB�~`w�>��&��(��R}þ�E����o�9�X m%�s+�F�����ڽ���%q`�y���S����9�$����i/F0U��g{���O=�٣�;�^a��SBR�pt�cݛ �d���[����ef9�KA�v
��\��|�̜$�JN��N~u|�k���\�6�d�/�1fTpxog�2���?���'0]��z_[hId�߯:K!\����%8����}|/��FV ��((�~��rV�ӓʏ�x1�A�ܪq�ַ��Ԕy����� J��R�eT��m�~�ǡl����D8��\ЃY���}����;9��}�rR�ܷRR	3ƒmͧ{��8� �(��*��XD��b��2K��z�
���ݵuK˃�)�Qî~ȩ�PNh���M�,)e4��+����gp�X.xtd"��U�gS�xmخ���%Ey����ۇ����ع�����)c@��r�?{�TlH���Fn�U8CFf���������!w��|#���(p�7�x�b��6�ii��}6����b��?tG��g�K�R3+�or� ?d�G^��2�e'}5��Yb���s��+�_������5��ܤDV9�P�ׯ����^�

��3��ׄ!Tφ@A{5�E]S_EP��GH�l��%��a�y� ��#���L��RT�-�X2$ز�L�ҧg��Z9m���D�\�J�+�rO�ijJ����I>-��y֕R��1�#��s��j�"�饻�FoP��9�*e�F��{}O&vd�ؖ���] ���<a�%'���FFJ|#(��\���-���XcU
�{m�.|�Fn��@���:`;��߂!�:�$��I��-����{�	�+BQ*%O{��N��d}��K	�����(��r�������}��`���6B'��rV�FYv�w-u��adх����ވ}F:&9"R?��@];�X���rb�SW��>��'h���Us��M6��i!Q��oS{9ʖ������?,rUPȴ_YK��Q�QZ�����ҽ��d�cc	2��]�ZZ*		�q��^�k#>�xlE'�
��TyN�����_�?[U�ЄL|�ܷ�����Рd��1C�^�J ��8�(#77��W��1�G�`"H�^os�>������_M}WW!�ӗ�֫���Q��1�Y�gUl9�_=$Z�,�XJ���Bh�>P7hM�$)~JF&=��(���`=���ֈN2��8:8`���_�v�xˁ���]RD�;;;�����bL8ʇ���^�N��[X�����d\�DaC#�:Ϝ����Z_��{t�w���I`u.@f�9J���Q�jk�?G[�܃�»�49]�����­��Nc��FCO�]��I A0�N;i<����KV6k�$��%�.�<���:��==������*��pGx\-�w��G��v�fE�#%2TTb�����7������A1M������ڊ�ܗPE���͈]?�'��B��hg_{ܓ67��V6��/߃\^��� >��zm�D9�̮]Y�3K������?f�f��9Ɠ��-��M~g���_5�l-#� 4���lA��ʸհdc�m2��h��"��ۛ�)�j������z)<�>'��)��K�anD	U�_A�g5�!8W �F	g���'MZM�vy��@���5"���9I�/0�;ux۬�.����A�N�*Ha��46�M��<90�QZ���_��k����y��mv
MoO��t��ׯ�+�˼?R���w7&&���\��}W��2�
�E
�I�Y���zC�Vq8�VO��z:III�+/��v���|y�}�.�2(u�٭[�~:L<�R��%��5����$�&�f d�@}����A�q���~��a"��b߬f�+K�U��S��t"��LU���Ch����2Y����:xP7�op��ܑ����?��k���$~6RH|(v3��7�~��s����0u��8D�T�M�Q=��7����}����ct��is����F�\��h�_xG�u�<07W&+�H 6�ZI9T�V[-��8��kO���"@��(�LN=���C3zCqPgHb�+)1�\�輏����}�>��v��0~ܚK
rzg��%%>�f7*2==�i�N�8\��5���?;M0���Wa�B�_u_M�/Xgm{�^]���<�<���ֻy��綩.�g-��R����oH����? � 4����j�I�l�����8���1����m�\T�q>�gk�01-1[����������z��%(����s^�d}�<=�����8`��XPK)��O�GEP�,�A���/��mis��;���k#=��E/�]lJMO�̮�0��m(�uA��:%���;��I��o=��0Fo����7��������� @�t��Vx�,��g&����<��.d���yVOSRn�Jk))�'�cHS�{�r����u��&[�{=���3WI��.�`D񵋬 p��'']��WM���kyz!n-|��E���^�sJ�X��.%���NP6�h-c�(���$mm�qY���ujj�е�������1f.i �[ix������N���1	�����v�w�c\GO���0̟w�)rߙ���W8�M�������:)�q��- �s ÈL��V�?J[��Ɛ-��蘘��'u�ZxV�1���c�Ų��t���3�e9�J��� ���*k�,���pt���:�
h#,|�v�r�[[3$qq�]��}��\�n����oԋ�pT�A�対��]�f�5A,&"�a`>S�!������x�!��w�uX�&�@vq��5sߠ=v|��� "l��q|_�[�?^�Tt�1fخ��K���Jyh�@$����<
��,|ji}�������F�`�^⯰��w������H�A1tt�+}c?V��Q?��'px7X�5ޕ�h�o��DN2~�8��2%%4��������f�A����i�!(��
u $��SR��tt|�����C�!�Z@/�o+�{�i���hbR&'�(
�e��қ�1�̋\S��$9#J���*�:��P�J�P��\�h��\�2�u�Jaa^lT�.�p�a�� )���f4����W��ǝ�� L���ό�z� ˤM`rI�?o�XWg��}����Ȕ���"��'�3��VT�kZzh�Ǟ�.ZP,�_��U�ЧOd2Y_�C���jh�f���z��!䏆�}�nI������P�#Z{(c���������b0�@�bv{go�8?��~DD�ݾ�Bx�,ϴS]\�_�M7�w)Bk�MV������=>	�����ק���6)�q����o�����v{�Lg'����Xk�
�����?�ne8��M�K�n��Dw&9"�LBK�2Bc1;�ާ���ʐ��3t0ם�B��n@e�**`�RS<�A<o��$�����1����W�I;��V�_�pp�((�ο{�A�w�6B&���ق���V�����*�Бf�]w���♹�0���V��f��jN��:�z��Ʉ�Z��m��l<���_���X�^���ʰ�o�Txl�Vj�-`���xg��ηe��8�����m]�@���6�_����Ԕ>lb���mH�hV[�44���Ԅ�)R�y���L7�܂��(�w�A��bP�T��b[*^dL��+烲��ꊠ���̟\���C�&&W��RdL��Í��0�F��uV]{9 �^V�~~-��E:�
Sz\]N�G3D}�,�jkڬ���Z�?qssu����0{j�(e.N�����a�`�+?���:�R��cN�����g���,~���FQ8�io%G����u9��F8�h9����е��Y�t��qպ
5��c5���S��oߐ�a��J'>�i��Q��jZ{�"&�j,����|�������@g�����K��%����$PZ��lE��Q��O��M�`�(�����11���}��4�V��0�x �s?jC~�E���*�@tԙާJX� Xu�:��=�:���΍��X&���s_nnL�R>�XB�,~�r��Iw-�����O$�6�h�ր��Q��F�皺�)�}�ߟ���������-Q?yr�P���X���51��Мm�u��#ynh�V�Ųk���c͆៌���4���x&��Dz0�G⳰��q��I]]�T��F%� (��N׷Dh�hB��<����h����\

�)OQ�s��������LK�ӣ��p/pL�&�U��V]�m�� ��a�� �S4M�[˓��4��8KT*�4g�U�=��s+&*�Ã-6Z����6mw��(����Oc��n��89y��'$AN��������7q���;��T� #��c����V�/ϟ3�3>h���Ş���#7�{+���_��� ,rjKv�wP8�_jjR��kI���K C���I��z��Z(��wuq�gap��G$-A�I��c���śx���@��׵u��Ζ�^%8)o�K�L��`�z"#O}��Go��)\�li�[�����Y
��Xik��JFn��--7�5����E��pt��]_w�Q�~NT�^)�w�'��؄K�� b��h��j]���͖0���=��Hv9���K6a��k�K����4�j��JKҪ,����eg����s�y�����Ѡ;�ɨ�'�z�i�x����0nϛ��b!�l���-m/�.���D��2CBs'X#�X��;���p�Ç����BIC�9kXY���˝z�M�JI�xQv��D����5�T�[IA�%:���B�l�A�F����A]!�zNR71���R�������z��*M�.O_��Ћ@��im5������h�jg�e
?6f�5�Ɓ�m��������}�$��#�r�Jˎk�]_~����WRD��g{��wvFs���㷁 �|��!mk��/���0Җ��q"��E��G�3�Jx8n�+��_�N�uaH�4��ڕi/�[0�T��&A�S� �0�GR2S�܂bKE�6�t�~=j�%P�90+Kek��tHH��"qyy�.n�K'��YpG�F�b"@ߊ߸y�#��{=�k,�']E�ȴPe���"�������h+�.���"q8�-�7n�fXXZ_��y"mHZ+�����L��vF�5g{�Q)�ʤK67?�%���%(9�i��?/�B������3���А
R��S��)#�����m�^\҅|9�X�{_�P[�ۉӒ��Z|�U5w=�1l|0;����/W�c>؞�-M����7*"n�M��h�T�1�,.r2r��/�X�Ud?*)��P��S��'  ����~��e4ZI�e�������h����sIL�5@1�y�p��6��l�;�K��ixu7���߉t�*,tbz,�D�d/]A�n��&Y��\��\��)G�e��Eʏ�2V��c[�U]�����ڭG-�,(ߺ�D}��,�"�2+�����BMM�x۱͗@oM�		�ٯ`�����-�IK;i25�_����;�(_��u�f�dѵB81u;������p�CY��9jN­wH��1 Z���|Z�O��@�L
��q��x(4����h�p���,"qgU���u ��9��h��~`g?�T[ۜ5�P��< ���/���d�*�u˿C���?��gW����^��q/����\9��HJG�;��ejlx�		0DF2X\�p��Z4�e��
��Ϯ�L�_bT4� �h�$��l9�X�*�B��И�
*�Е�į�8�fnvvН�Cz�-=lI$���dm����{�e��M�
�M#f�k��X��p�z�x/�u.8g�
�����AIO!)��T�č�Zff��y'��܁D'�x⋲���iQZ^u����������sq�	�Ѕ�v|�wr���M0r;�(��}�����z�:K|Hp%k�[� �;q�|�1�>.]\�$4t|תʲַBSh�vXL���b��Ћ���\ˊJ<��
M�ſ-����>��3	ڞϩne&�������i>ܛ$>CfP��d�_��Q���Z@�s�?�����Dc*F�[k�.\�{hx7���u��:�l�+����i0�qK���(���v�3�4W���N�I
�M����]]�=�M��"�`ՙ���b<^�86F���j�*��r�N�Ec^;�����(���Տ]����<�#Ǒ��;���n�&2j��V�5gKc��Á�(̇�[t���T7���2F`.d�/���ė�O�a�	1j��>�L�}s6�mss��F|����i���Q��1r�( >����g��鍉/�'.�;T������2`ND��)�(�eF~(4T��L/?YHIq��p�6Y'W��$�{]���ϯ��`�#G�Ǎx���2�m��!��~�9�r��҆�թ�MFɬ/P�i�����bԨ Uj**�����_u}��ыJ����>F�4{�)9}��P����4����ќ:�����X#�]1�CR�wa�UW�-z;3����|"i@_��DI���Xr��B��U�B��.����;�z�;��A~�ݷK��%i�6���T8�����:X��x�=��4�i��Q?�Bݬ|�>�@��h���֭3ۆ�/�i�ߦ�_�>hR�H��'>�W��XK˛k�ܮ��ZZ����������X�5��2�k�vq�$b�e�"Ū��l��PUG{c��l�k�Cӊ {� ��n�4J(*L�vu;�^�G���Zd�" 8.9x��V���FD�C-���j�C�@&��l��J�M*+5��k�9�i�.�e<�!QQe��;C�h}ԉX^/�E��ep��E)��G~�j�n��j6�����O}̎��San�q����O�$�
(o6#.zz�����bNX��[���M�l�ll�@���s|i|ӑ
E<kKZS�M��ׄ��<36�[�O \�Lf�X�h����_C�_���X&��,��ǒ�.�FƛOa���a�{�OU1/���7�@{x�OSAM�Q��w`�����5�k�AA�J������>!�4�qF7��$� ���t
Ž����)�_�� �܃+k�q�='��R4�kr���	^m��[5�,
�|��3/��#�E��wI8表~��1���.�(�'67���
�}v+#�J��S��Ђ��0��z����T��g	�\��?���{��x;��V@g*��1���`�dC��k3�J���CG�$a�'�Z]�����Eig��P�>JRP~������.��QM���|��fa@��Ȼ>^Y�6����� a�&'�����[���p[��"�Q�7+{�ui�kC�|6袵��Lm1��P�⶗e섆׸Y%��* !_D0���/�oZZ� ��]N���Jq�e�Ǹ�k����Zi��b|���:;-/�O����������]�^����DA��?�V�����d~~q���¢�t;R�-�`��%y����QH���.�qʌ���6�鋵.3EG%^��c���$������O%$,^�1�!
�T"x/ܟ��ΞYT����; '��hJ���#%�8�]@�G�j0��82�+%2��U����h�˴�@>L�lĠ��m�0��T���B�}�6�ݕ��@����ԙ�k���m!r2$��������k��0:L�B�����A&`t��sV���l7 .�_��*��"I�+M���N����&j~��ϫ+CT	V�����F	BN	�@8��S0N��)���<�h?	`��[ b@x�>,����_=���	v�1x��e&���k�}�_Y^�b p�*�g}l����y������,@zl�9p���D�'&�$�&	;�gxه����:��NWAD^��!��wMG�Ga���̇�x2��K��X�f�� "ˣ ii��[�-O�M,pB�e��F+ˋ���Ê
�����P$5��N�v�U:U�['�}ț@��e�����+\Ζ��wL><j��A����tt�A �<��<��6��a#}�۬�3(�-+�ҷ������kkׄ��)�O�lA��NMk&�͓\���L%H��k���=9��u��O]YQH��ڠ��d=�%b�a��r8��(�N2<u�\n��J�{���� ���`W�Mn![:<��^�IlW��w`�'��ޏf�wu�^�g�0�w���(�3:���p�iy07�	��Z5CO+��^C��("�7������DS�:	�Q�Z=n���$l����E0�(lʰ�44����P���-k|�v/ņ��Z��)��Cl���f	�!:-ϒ�}ך�����m��M.�׀vJ���V� �g��������O��I�t��cq��\�fIHI�q�����-I�c�#��4�4v@�_�+*��A'z���fK<�k�a�{.)�N.�0S��1iP������@��<��Z��u"�pӧXX'Z�e���,$�]q�L�Rݥ�V�u��[7[`I�\i}��#��$FF2��\���K�`����N��xp*.*��w7����?}"]�0��X8�+�{�t�<{�,F�t`��l]Mʳ��?��Dm������M�<�
֮h�<��>���_R$G;}<�َ�ш~M'���}���}yAi�,׊FBw�I�̣��e��O
��VL�m��Q�����'-~dS�N��t��uOο
��j���r!�	���t'�7�}N]�GU�����o�7��mnZ�W�����2���3���%���ʭ[��s����L@�h�)��͌��[�>�O^�1�!��AI`�9!��d _�[��V�s��_'ײp`,gc�礯/,�kğ7d�=�%���OC�K�����蕾�$���w��sUnѰ�{�S�)ނ}�x����8j��|�;���a,)�m�m����I)�=1X��N��������%�=�5�<�B'�b𣞫 �*����H�
6l���G����#��8�Y�x��h���9MQ�Q �D'�Q�~R��?�ctW�b^v }	k�9����Çɾ���{J���A'�G������|J�y'w������W�_贮��(h����`g	)(��.���
ߏ�Y[.�v�����	��~4���$%K��ߡ���y�,
�k�/�ΩU��ԍ���-�MA��gB�U ��*���
�Z[�$����*z�	���g��������@d!�s:�9J�Xٛ�����R#�S"@S���E_�n��+��NH\Gt3���z��ʧL��r��q�Qt� zj�u�=�:�&�6|��f�J�֑��(��{��PuM�w�ѯ2�(��8s�W�py��	�$	�ߴ>��Z�b��Ǹ��*@z<*�����rr����x�^7t��<��Q�}�/��)��o����]�q[�7Wl�����Z/{
���F��{��[_J��>  �#�N�%$����C�#��*JI5�/�w�K³���;	��mp~��#H�If�꿠���P���|��4�TUf�'@�T�mI�3|���(��Gu�������4Y��7�����&0H'�n����H�]Mqz��,
���Q�IuQ��@,�C,V�e��W���JȾTT=�b��@� �FQ�};�����Zd������Kqv��-L��$}�w���2V��_���4/{�aRC��xYZ��X�%�q����J�ͳ�!1GM���K�*F��I��;Y���2�i)N"����둯9`�g�݃/-f{�T�}�����hj��U)Wע�JK�lN��ᗾ5m��A�)x+�#[ڏ�����#���5٠'�����_�9Վ3>x����O`()5X^��t�g~E=��s��l��p[�"y��Hk�4������B�]�0R�}$~|L��  ���~�~����4w�)�Xָ=�Va�!�^^��#���}дG`.ɔ0zlu���ǿ('�m���3m����D���f1�7?t�T� ��i/M Q�ꞝu-h� �Z���\�,��a��M����u�8��i�pt���Xt�ũ�J��5�nA~s�:+�_f��!���l��� �Y�I�\���.�,�z�ɪ�����o��d��;2´"�ߌ%P��{���IlR�!���<k:8���XE����4�~!]�g���5��yd�L%�����-��]��w�{��(g��_2�U�e���E����~t�קaa�}Z��/2����v�W�g�Pńw��x�{X��Tw�{�@�U3_%]���$�j���9���_a���\�UAM��ў�!h�O��1�"�C�g��|=�{/	s%O��/�U���������XŤ=�����.���4�4�VR-���h�%� ��+˜�&��;��^�Wx�L>�e��Q�5<vH�fB,] �����;t�a<���P�R�*��z���C�(^��89���8�(B[�	?�C�zY�o
��=/c�"t�?�t�+[����ɲ���>�2��|��I��r��;N��{(}���|м�0yeC����n�%h7�!�dkLn!�%N�Z�	aL��,���EB��Wmu'䒄�Sx��M]>��g�g�NN����� P��������ꊕ���ԏ��H-�����fろL��E�=΍���p'�i�H�VR�������T��'wsN��7���٧�DA��%�������@Cq"��İ�YQ���� �=ݙ�e[�Ԩ�7]ب(ttQ�nH��LJޟu���Xzf�~@0��.��I?Z�}��ӭ!��Β#B����޵�t	�j��Bt��>�W�����Ԓp6�x�8�Z3����7H�\��c.�&J����,�Qh겳׮�D,v���u�O�$�6�����$z����={v��*��א��	h��$�w�f �t��,��_����ٍp�ٟc�K��L��0vp��T�. N+���m�]�{� ���m�'���q�h^�.:��/F�k�!_9�)"�I���H�J��ϟ_2�:l����o� �/^��^i���;1�j�>�=��6�K�Dr�.$0>m���;�	,6��<2;??�Ț�!���׷�͸�o�����;l������x�����㳝#�\ۏ��S�����^��R��>�L�nj��#ܜ�:�?-h-���)a��v&\���K[ŞJ���O���xɀ%�Z��?���cw�X�|�4��O�4�vh:��EUS
�zϵ����
4�{�X����������� @�S�`�)Ǹh&�z�.�����O��Ӝ`�l�FL���i2�Ny���y��F�21��Z{׌��㨕�Ќ�i��˵�ҙ�".���e��E�(�]\��@��+ ��\�T�RxKk�+�#�dZ�+k�<}���p���%)t�)���P��g|��#���	���ieg���O�+�`&�[k�*)�Vgd�k���w��|~OD�w��5��n����5�OP6 N~#���K�(���3���/R���.k�juI"����8Y��.��C�ss�����ș��2�J��	.�a|��;#B��m����B���dL��u<6�wK�z�yHē�*�&��L�����~o=y͕ܸ������x��~�Z`�Pp�o%��V��%�~8�Нm�[4\h-��kp�*�9���ص60�����闱��G8�aDD %�[���Z���(Ι���s>��y��+�.�����(q˯��oEv��d�]��(w/���{��{>��9�+@��tgK�9mX��ɞ�e��ޟ�/�{�O��|v��q��Y�9��nm�\~�{"���)"���|nO>?<��vz�����*�M�z��X�ޏs�݊�ޠ���@��gy��I8Ԥ�*_Z��Nl��y𜻢��g��Hj�(7C��x���&p�b�M�no�i&�Qi[�g@�/��0+8�qh��dٚ70�~~���p��+]����]�>�,	�\++�Rj���Yߞ�c�4���n�����f�8׶H��������Kw�.gYVWq��<2p��3��^v��K<�����|���C0�{$NZ_���$Tq���{I�@����ڬ���%/��@k��&j0�ss����5h5�ݴ��Ao�͹�ϙbQ�Jt��wF\�b��7��DӅ�!��`�R�fg�m���>��+����a፝��̸d����;�a��K>̅V�����ӣ2MT*�{	Y�����Y	��W���@<�cC���[ݎ��V��w�;���9b��
�E�%i��/��s��i�~oRW3�+�[�ML2�w���{���#̖��д���д=ר� �E��NDu�sV���ϪF�)~�_w��>����nH��>:&I@�$FG�UuC|��!J0���@����GS�o.\�鿨�h�Tij��{��F_���+BA���2��}!��U3��2}���_&�^�.:R��;9���i��L ��=;%e}�n�K*�{�ueŝ��΃e�:�ϕ��ؔi���d{{{U�77��@�'��{�B��ZU��Z��T�*iE����B���{Qt�l�]-L\�R?�a��<?�ɾ�b��s>����~`n�2_���-����y�(ߔ���6I�Ͷ"�i�+.qpH���A�!d�U� 1q�ư����qO`ڛ���B�9�z������N���[���/7�+���иDv�!e� �|�x���+�j��_g�̸z�;���xn6�@W��^�@�Add�a�u�"���2⿸n��!�%�c�0����,�]���^�T�I�T�`֏���)�\��@z싈L��6=�-��H�<wmm]�-�����O���x��֖薨��'XAԻ����-��'�s/��<�dC裹g�g�v��'�
Y22/�ڻ�<=�
��J?7�����w~k%O��77�Y��y�S��ŵ|�{��g��9�WQ1@!���}����"7\\�������CsN�CsJ�w�H�&;@v��J��x �1%dc[l�2��g�Nb�&�!��2�#&t���R���V�'�ÎC��v��� �U��Q�Q�뇱�����}N8�����¨(��?�L��J{��dS����F�^�+XbH5S��R��V�H^bJ�Y��/�a\ŧ�l�A�\�w�	�P��z�O�A,�K1����2���F"H4��.�D!�5r��,'�}X~W�ʜ7�r����ωJv�Ƣã��y&�Q��g���ggA��
 ����I6%v=Bpm$h(�~F��"pc��ɧ����VB�=���y�4R�d&#~�"UX�8�ʃ8a�&�T�ʺ}�</x!ax�,��-���@�YTb9�t���U ���;�����r	�^DIADE:E�KP��[)��V��ne�ai�.�����g����8<��33�}�=��y�O�|��,�k'	���P�T���{f���ec�{�ʏHD��*�/��X\��uH�%���ү^���Yȕ;��G�3��R���j�=sPr�B�]�{泛S����
��<+�$�����^���F���O��4�Ź�&C�\1���с����Ξ�O��m+Xl�����(�:��ڝ�GW���.Pvo��yR��p5'��:b�_Y�@O*p��Du��Nt1��"ՙXP���f�'��p�bvy��EF�D�*����w�?����!Z����!�̽�e5�h�z���&T�]���R��ThLR�9�X 7�����l�����NC/nq�i!�u�O,K�K�+�urf��vk81�ʄO־���#�Q��ږ��9�u�0�X�s�]NW�y���U�p���rIx%�b�	�\�B`� �E��ilS���H��Lޤ]<����h)�kf��?���<�e:@��U�紜���u��:�����7ׇ����.	��?^�r������c�G�۳Y�[��Im	j�c�Mv_���k��iV�HP����v����_�:Z�';�����L��=�C�v,�D�`�����`.�PR�h)+IzY#��p���|ՙ/�1`�bl���՞��rX��<
�xJ���וH�r9�@
�9��Z��-�X��6���i��mP���Ik�D}�]�onu��AU�X���^��S`�{R�n��<�澁��R�7a}���~�+a��k��!�v��1*_�vKn�T��>d7���Tn�}sbA,�%yj��T�!�`sݖ.c��nL2t�w`ʢ/�F��#f8,A����n���=j��z(.��v���:�J�͆rqm�V�� R�;6���他�
��Գ�_�����v�N�\
���$�[��h��";���[V]>?�����1�J�N�?��/G�+��2��`��vw�+*":������w8�y2����zh]'�nWex�Ӂ�s�o��"�-A�%�jC���
]�x:D�2ER��^;�Y%������Y�8)w�ʷ w1=�W�������W7�b��`��Wx�b�vw��_����$�V�*�=H���>dp�3n^ǎ��������xNg֍]Ѩ6,��G=��XM�g�|�@R`�&�#�������*|i��%��P1��P:�0�̧�VC8d}_����%w/o.�}��6�\��"h:X=�_B�6�4#H�b��x֡�!��$�p=S�<�QC�А\��>翻 ��R^�sv�A��{��C����c����R;�����Nj�&̐wpwޙ+���o{�5��$�e��:��qK�9o�8�L�'_rC�|?teJ=1R}[�\�QE�f�7?�j9���V���AJ�ȝ�Ro�T`]��D[�uĖ��Ỹ�����(uv�7�'��-�w[Ìg�*��L��A~�L23#p�����ٛ�:�$!#�Q�t���f>�P�ce���:n�R��uH�Ҩi�M#-�)?�_a���3>��r�.����$�н���3�y��F��$p+]Q:E��	�_��6�^h2Y������B��
�f��S�O=��%�v��T�.�����l,�'������M0�͕n�^�&pX���[ ��
�eʿ�`%���ҥxJ3u�֏���+�R�I\�߆2�bѹqDn�܃G��~����S�p��#���jSH��>N .T��+������~��?�U���Zæ�X��HI"`-�?ɐ��XHov��i�"���AoT����UЩĬcUSw�+Y ��q���eN�� )E2R{���ϟ���gu�_��\h~�(��(n/<�:��Q}����� oԕ���^iW�_���)��S���=�>A SR��ʼO�r�0�?���+ʚ��ߺJ��n7�oq <+PU�P�,cN%b,�*��\�8��ܜ!_��l�µ������<��;�l�����c��_���V��y:�$�^�ٟ���`�(?�n����9>9��6����k@A�SjkJKk��\�MsYX&c �&�+�Rb3S����ŭ�}W@�g����R�#�����	4��87��W�8�i�"�.�ꁇ���V�����-U�>XP���/)9c��x���U�:��r/�>�}ZU�v����h�Z���a`��Z��Y卺���c�W����acK��Xp����6�Ԕ����n�H��U�',>��7�nni�i7s)�ھ=pK�Ǯ�x�wdm��~v�}j@y�����cƨ���NsC�껼�D0�sڕ�V���}��b�)�[�L�])�FH2�w����2MȪ��>|W�� h)�h�?ɬ�c�
K׿	S�G�bAA�4�@Vf��.s�^��w��C=O�<t.M����9�-��fG##E�����V��V��-zn5f����MZeE���d������X�]���l�H�+�$|q+�Y�!oS5�GE�yr��x����G�kD/����M��yv{j�uu}�;�&e}R㒦���lf��=\{�g;U2����M*�.ì-�_�%#����u/N���6ܘ��!�	`=��>���?�(rm�j=g� |o�
sq��\@ѨUځ�1|7�����O�]�bN�?�Z���,�T�$a+JQ��{D�Sw�b{Np�D[be������^<�ff�}^wE�_!2�$JKH>V.<���݁�'����� ���0WP<�xo��U�9V�l !��j�VE�����	�:�~JV���a���8s��_�|�tg~f�1%�.�θ\<f��r��B�#�_�`_���*��7F�#JJ"�"?IJ�&��zIAu�Vz`����yHXϔ[�A��ʕ�=���K���hA�"�2$����mO��]V��[�y,����~1Xvp��ZJO���P�I�j�?՛���~���qh0�]�vv�=7u���j��=�T��{:UfffeT}_]�:�HV����:�d��t�>���\A��I��	�xn�6��{��>I:Ï/��i��h��!�����6�#��w!_���8ި��,E��:��'n���
��k��-�3��9%�AJ^��,--��x9�i�1DcՐJ9Y�g�6���콳p����My"����p��v����ڵ�]�R'�E�s�у�3�jχd�/�ʒ	!�㉝jz5$İ��j��E}֟�󊮲3Q�k~�]6X��1�������lyg^hE`vN	�K,S(5�&Z`��p��k�����,Ht�颣��	�%�A�n�ey�\R�����s[��d�7M$/�9���qN��r�}������T�6������5��L��R����&`$�e��GP����И�:�kH�W�v���W���\�°�ܯ��q8-<e�_�"���ú�~_�������ڠ%����S���K������N�����n �������:_1��*�t�_�O��˟a�myn7�\|��@�$ �	
���4��9�Y�������acl�z闱��BC{�):z�_��Z\����șt���W��y�ya� t����#�|���R�4�]�҇^�O��g�ӽ^��`��"�AqK�U�T�຦��M�&��jF��c�}�6�g��u�~{C�'!!�b��?��� S\Hn ���K��]AFy�O{O��13��/x�~y�- d��+��<N�e�O2!Jܕ0�s��S����8�?���W�������~<��n����9c �4�J���q����p�)}���oyi�.�;b6p<���Og�9Z�O	B���>��֓3Ǳ	�
��|{�x�.���J�	��|�>=zqUf�Di��s������y������P�����Bd��nD([��x�)��γsx�R�*����BՍuT�\�^$�O}��"J�0 ��,x*Ͱ�������m������/�MG����cy�M[��J�Q.{+�-t��/ar�[����V+��"��L�e[2��h��
cVr���TY0�D=��Q�3ߚ����M��P�{�:l\ 7u$�V�����~70��Gs�W4o=qj���y����7����f�����1b��D���XTbd�T˩��Y0�[\��tB����C/�`��)�_�'0��d1%���I� �y�|��ı�EX�,�+��H�vu�=�7�rƑ�ii��y9Q5N�s���:�v�L�n ��7����4�f��(CƧ����v��i?�#�����Iۅ[(��9^[�_<� �{p��2�v�d�{��|�)�)����1��$Q�2rEV����@�C^G˷,\��]y(��m�����,�Wb�����w��ff^C�C�Fs�2d�F�
^$�\�++�Zδ<2@]����\2��0��¨+�Pj����F#4������*�ǃT���P1M5��>��eQwF#�]�P`��w0\�̬�&Es �O�������.��*j[p����������D�l�l5���R������4�D�ܲ�Ng�t`����/����<����ꥊ��;,D��������!J>�4����}�s�r�����l�;o2�MM�JA�ƉWe>O�H����-�1]���j�k�[3�ƽOGmq�#օ�2��+����ػ��СV�d"�������$O��@���V9�0 ;B�11	�f����ZWG��LE`a)��1�(}|܇����C��o�뫬���Q�p�/X� )��n�\�(Ri��:�=����f�~-�	�[j�Se�$��{WY�����ʻ�������z�v��`e���m7ƿڵ�.vx=�1L�r��@����vK�z$c!]*\�ݸ�j���щ."�ә�%�d�EQ�c���\n�W���j7$0�'$�~r�E�N**E����?aT?{�ۖ�,=ѝ+���ji���]?'������L���~��m�e0�����:�������� ͆����}'!]%:rM@�8j?R>����m$��~��4T�`�f����촄_�Y&�jj0�r�s��)UB�'5UKk>��iT/Z��>��1G�%Zq������!7~Y*dr�v<�%�	��O�wR�6�}��t,3��H��ٵ��УNH�zc�1��~�-30��[K����D�K�Y����c�)�Ƴ��iN�t\�&��B��K:(��������M�|,�_��3MDw?WK?�r>	�l�[�|h3mtL���v7�rѱ��0J�'7�hՌ���yd��2��[�}��*>���?Cg�Fg��{	
��Xo�#"��AR<�/7W*������j��� �3�)�~j�<X����)st��}��?O��N�Q{���`pi"����@M���/���آ��r+y�� �'n88��8������{tq�Q�L��`@�q��w>vf1wµSR������i�́��^����+1 !����U�k2J�V��� ����F�
�Ry�;Y�O11��v�_p%̿��*b\�;��A2KlSIme��6�������V�"�����+6��u�ȫ�Ulum0�'ǽ"��SS�~��)�r1�U�K~qd�˺���i��P=;Zp�x'&
~u�n���&|�
����QYw��7?�bLZ�[���Z��k�U���ANU���7?uV�t�?׾�؛�\U��£�Bub0}5������{Չ17W#�$��ibl�(���h7���1+�ۈ Z������c���?0�;!��6<�uu� ���Ɛ�GH����&��B�1ܟ�S���|�i˪v�x��6����	��dn軉sS��0�N�}�ÅI�,�,���b����i�!���� =�l�g
`�|ߋ���'���N+=ۋ�%�M�0(�M8m��4+�g�!%���N����i)7��Bk�h�W�n7�����jq�����+$�1��hL�����K}� �eU�!�Rp��6i(h����_��s��
t"2(J��������C�z��Ps�߰+}�wAJ'h16v<�n��Qا+�2�b��s����_���?sD�$dO���M�ڝ1����b�R�s�ׇ�%�.³Aj���W����X���V�7���#��]ó�h1팒s���x��W�\��8���pMM�ט�@ʄ���'��F��!��=X�@W#�\*�[z�iC��{��4�I���?b:�w�/n�!eE9��{����3����E�b�H��`-�+[^��Aly���չ�Fͱ�>�YJ-���(��F%��/:�dp��>�/ ��x+C�^i	���q]I"�9�B@?,�b�{����Xl���h���B���i�;b&����Y�J(+t�!����Q��J�Lzv%����Q��F ��]���$;(BO�Ř�q���yJ���FY~ ��T��s6�â��o�i7�f@~<[���c�>fwu�5��`�
��7�$���%;32*��DCuL^Du!Q�y�C*��W����P�E$����W[@�H�G(o��~����������	L���P0��b`��tH���]NG*ͨ)�^ڌ�����jH�A��z^�xu��&�aK������#�Q���Kx(�	k���x�u���T]'�v=��Z��=�DH2�����ю!��\6�}�Y��gDM��,�5^_w儾���d*�ۡ71��[���F�+��>��2��1z�V�.�'�t�2���,YԵ��BT�ʾ���f�?;Y]�^�-6]��p�'��Ƶ*8}T�����݄ZqSdi'N� Fql�i^��::Fʑ�}��t�{w����եW-�������nNz����G׀Y�,/+�n��e4�!?�eB]���Gi��4-��e�����3�~}�!��R����MM˂Yh�δOmIr�����-'1��
'��>��9�n��$nnjcMҿ�,�1:�
E�Ʀ�g���)r�\�����ec�j��n
((*�]���ϳ����G���9��,/�����j�t�j�rt������ͬ!�؊P��6�`G�gᣓ�P��Ĵ�y�'A��G(uqޖ���V��%9�2]�=��k��bu�5A�{H�]gwp������7�!#Tw�m;]<�� #D�Y�tB`J�6y�ܟx*.frd�Re���j֑޼6�]1}��3b��C��(/��ܼ�i���>їH�|$��yfq|�'��M�.��,�_fNM���?"$6R}
��9.��@\��=?����2�Fs;Pmj�023H�tv��`�}�������=���Ѽ�#�d��
2��ݾǏ�����?�M��s�!��bFjB�\��O�J�r�񣝣	�TDLfU	 R�r;I	]��t��F����_��n43#pp���<ݛ��BÅ���s�0	�\h�����~�L�LKН�^9y���'�gw���O�6� ��P�=��!Y���
t��9 #�}��s6G-�硰(&^ݫ|��{�sQ;�??�iv��귯��jT�{�����d�ٴ� 3������*�,������)C��kdEG��2$0:Y��\Kh}�a�3���5e�u<\�}�-�#%��)�1���M���Ѩ)ٛ%��"�Aj�~�0����۾�K�ٺ FH!}�`T�����T���L�9�G��|㪛��Bc��EF���|�I�\9����Go'O/;?u�7��>�#����� �D�������"G�B\X��:UK�����DU���_G�n5 �%��SqJ9�tb_ϙ?�����j���u�yX���gCE���M�:�;ɫK҆�ӹp�`��Ų�.��zL�? `�E��~�]���}�g��L7�i���JO'V�ȟ�-�L��h$rKCS��2kԡ�=d0���A����ht�J3j�~<��}�^Q��6�РP��yy����du:��BQ�">q�c%��Sn�t3�n
�@����Ё�z�T�""G
���dyu��I�:�Zna��c�a�b��I�2R�g�Ǩb��\\�ڳ���kS+�1٣���(��.�H����b�v����>u��ϝf���7Ǥ�p�<�BG!���M<�vO��NIɰ<mi��8����}�������W>�u��#3k!��3
�MZ�΀����8���<�a�Td��r 쭿uBr�!��奬�X�m����&�z�����&j�8����A����Ŗ���ezŬZ�}J�twG)����D���ҐŲ� �u+������̼������w%��| �b�	2<s:��D e���p
��5eܘ����!Jƕ�w���͗�>�U@��o��/4A�o2n�|y���P�6����0�z�����8�EeQx�P<1��~����[�g��b����a9�$j�n�ru-��=y��=��5Zu!�	7ξ�7�i��c���!DI�2�X�K�!�][s��w9ZT�(�ى�|�N#"/�2@�a�����P�Ú�Q+��it8Q��;R�#WN��Z�'�)� �	��B^M��O�vg�nIJ�h�Ҏ��#�	�7�]��?�q˚��q�5�!::��I��%srl}�����5h��0h���"���us@�*]"J�si�n��n�oM����u`
Sj'���f�~��h�q+��i�ٹ��l<�X,G�����u=��Jz��1���p��Rɏe#r�f��6��C���I�de=�v�2��U�E�������8�>�@0�-�b4Szo����Z���M0���_�Y4���ai47/M��T�cb���{o��#��D��guL�rۉ�YBDީ E�!P!'.�O�u�^�XLy*`x{R���?:��ۼ��7���1)RP��|(J_��Д[�kux�����tEEE���c@�<>�V2�+H��r����S�����ǒ�W�>�	_v3����+s�Ю�ANŝ眸a�)p*��H.v ���1�I���En�3�
�I������Oo�b�t�u<��\rW����0��V&����pd���[�ۨ��eSa��I��mU|�N7��!D��S��D�ff�,|]:P-� �ws�CR��lT���M��p���u���}��U��ڋ���3��D�������bP09M'Q�V�`�.~͆��'ׅ���B���^�U��(�8�}�3/�n�ʿ�!_Y��:����P�<��W�^��z����7�4���p�GU����	uvu�H=�H=��zbS���$ڶ�:7�é�Ԭ���آ�_�=���1n0ra��d4��z��F�"!.h�I�Χ������6�F݉�.vZ��<-B�{��'�Į���&;0��YoX��n��){��Jt���g�H;�W��@m�<m�R=8OS[�\Z�ȵ�,��j�g�c�O)�1ZS%7�+�>Q�˂p���ӳfoH����AA�xL�<,�m���.�B^�i��1ϒs��kOy�<�!._~8-����-gv���=u=L�~{i)�q)��F�����gVK��K~w�ܷӥ�-3������7�R���E~@~��g�y��N۾���B���<b6��,"�bk�'�C3�B�AY:>�#��w�Q�و�P�B�_4��qX?c7ư�)o��U|���|	��o���V�Z2�h<�?���U�D��o�va��?y�7P��_����W�x�^���q�װ� �:�֬��u��Nb&D��|�%�]�r�oENR9;��ȏ��߹�8�������1�,���	�{�oLy��|���Eb�Ϋn��%f'Sm�*O~_%���^DYu��Xy�)XHz���Aj~�(�h�q����~����0�v����2<xx|T���,!��)1�g�w\�L�G_G��`"`��[���*��h<"l�2j��pГ"=nNBt��>���SX>ɘQ.�U��HR������ގ�l���M��n����uԄ�b�� d�z��Sox�[~p=��*�0��z g��K�����/Ưr֐�_��a��_�)B	�-|�tq���i�����W��Xd[�Gw?���6*h�z��x4�(�݉g[���=duGr*U�?V�6>6�L�ݒ�����_ۣa���	X��n����V�̊R��l�5�+.c⿜6@�����ƙ��;��yC�^�-x��VC��WI�n˹��5%�\8E�V�?K=.��埏��>���$�� �ԛ������r�o�u[q5����O?���DM~�8�۴���=Q�,�u�$�{��H�i�:�9�����Tkn+�B�D:S��ϖ�ͺ�5
z>�W�E|���^�H�VK���1VFRϛQ]�*���-C�PX�^s�����B�t���iːV���;7^�6Dbt����/����#�Z*)b(�(�!H&nn.P��w�×�x����xSS�`�%�RS���I��P��оJ;���2��c�������E�+-���P֨��0�e�1�r��̮�^q��Œ{���_^���\;o�5����4�
rΈD�^<�j�V���[`�����җ鍍|u�t(�P���C�$g��q�k�qQ�)�`���G[��[��B�M^�Pp�DFy�{�����>�0�E������z�gޯL\���2�V˪���x���NK����S EQq����$�[<[X�m��tk�a6j,G�����S���b9Y\Ћ&�:��;kW�d5�;}��#%��,M��mr���11C����7[�/X/w���G���O��]�u�GX���W��:땓%��-��;9O�yAZ��#ڠ�@���8 ���q����Q�rλ�O8��Ū�v�+�2'�&u�pQ?�2]G�4%�*���>u_h�a�k��p�Ͱng,�5Lo>��x���ShS����;�D�l%�؉g�)o"��*횳G;��_cM٦qJ��mp;�	A����}KLO�m/�����3�*79�
�jN�q�e����e���mw��	 ��ef϶����p�׬wd-��C�����Nl<�Ȥ[����� �"N��	.G�pt��%şf���)H��ĸ�"7W`Q -�C.vH����q@]�x�jd�!��� s��9Z��F�پ�Q;Q�W�Q�̋���3h�5XcY�`ڝ�MA���Dc��dl�^���*����"�A;���iFT�G����N�]Y��)�Q9,�4�����4>�y��g�on�vN\��C2sN���"��$����������J�j&Hm+7�L(I\)_t�}(Ğ�Xf��T��j�UW�o�9��S������GGY��r�ŝK�5c+G���'-�J��J^���}�J�i��Li��!K6.�����T@Hb�#�K-�)�~68(s����6B�F˼�UJ.s�V��[�Y�B�N9Yd|���<��Ȭ�#F��{���qv ����"�dGs�0���>���i	'.xo75���aA�ؠ������v{�岽I���M�%7��iT�9�}�snX�h�7(���ѵꝦ�	ӿ��{$cŔˋ���r�����I�U!�mc�
�G��A,�?zR�/_����@�#z�^e�."�n��i:LG�����A�a�����\�{+'���?��nZo��VI��9Y,B7���@EG���v@P?"��Ŵz`��J#�T@��~-WįE�H�9����F�m��Z�R�����J7^����;"r��A���.R�@	�C�1ж����mm�\X�g΁��,q���-»\��/M�
�F�����9i���$���x��ML�(<�k�dC[n^6�Y�~���t���9CT�T��:�V6҆&(mdt� ���m���!�G���4�%8�� ��̓�?�V/+6����Z	�o����w;�[;ItݖB��aPQV�-AI���� �����n5�s>�^9��.��5��@+�,�L���Ifo�b�j��ˌ���+�����OI��;Vbb�]�q����K:&S��Ϲ;0u��3��-d%}��E���� � ʶ�yq�'#)�f4���  ��θ���,�����֋�P'��Q�v���"��KpqB#e���14T����̴��#�5��*�Pv�����i��a�a� ��gb�
�\��S�o�1���� ���w���m�iv�Y$K��&-�;b�</��fВ�R�d�p���o�o�b��E�>r��4PY�L�#�g����S�z�?{X8^��B�[�Q4��TZ    �֕�7�������G9!(�(���ZP��G�a�+^����r੿6�9�O��V���n�
��K����dBU>*���s���9Y|��!�)|4�AbΒ�1���j����w1�7��r�-pO,��7�+���ȣ��[	@��'o����fB�ŕ��x�I,��� �u�nA����DS�`%P�
9���x��d��ø*s��.���V���YɃ�)�E���{�E�JY���*�||'��N��R����"�;��YG�l<�Rt��mHS9g�^�,�a��b`���=\���ѯ�tB�w�O��Khh��~L��uy���� �,ʉ�JYq��
�y��m_�~��v�]OĎ��������� h���娼�ҁ��J�6�
�(��&����`*��<ˏ���LJ�-���{8�h����i�T��M�9�F/����Ncz�k&�b� 1I����y ki,-�p������x��L�@_xT�<���>�pM#rif��m�,�lǂ�����~���:.�YϺ#�� ���]kF𣰐�**��Q�Z��vʼ���u�D����^��n�����b�y�d���M�l�Ҩ^-�w�e�(�x~���pg���Y�G�8[3_���]��`���Nօ�>L��Hgݮ�p��Ąہ-����әRͮ��T�p� 2�:��P�Q�/3���~T�߰��^E#����<��@h�dQ�ו����	|uhzx��<��r�w?K���'O�Δ;w���~��!G�����uU0���?m,���(,?Q[
dܷ���qӖ nTt�<?�$о?V���(��P]9{}ܬ������נ���N�.�\Ov���Ǿs3\��ڸ�~ �iA�1�G����X�I��&��A�m�ϡ��-��Lq%�i�+��3e=NFI�*V�Y�7�O<9"�ac���1�L�)w�M^&�.eX �Дկ����j�����DD�SO`D5������%`��Q�j�I?����`�$��`�� �n�wet�����(��K[7<���n_11��!�%}��b3�PGqӏM�[h?�ɐU�[����b�15^\�u0J�U�V�����}�yA���	�K
Uj�>W�;K� U�܆�-�'�x%@׉HOײ�U�8��jm�8�[gLdt�h9='!���]!�P��]U6��H��j�f+�JLǛV���U��8�:�1�M�4%t��%t-<�;m�t��h*�|��=(�K�'���i*Aǌ�8�EF�;��� �8܀%�&�Wr�L~~�V!��R�B%2Q/r��dnC�k@�U�RwWב�󍍘`�sT����Q�o��,�����\��w�,&Q��Ѷ��Ƹ��&6B91����P���<t�y^���uT'����0���4��p��i���`Z̔9 \V��9Pԯ���6޴T�<ݖ'l��$��d��2��RS.��E�1��)B�7�#캊�7/`]~ ;A�Y� v	��Dpo�����*Ɔ�8g�����M��n?r?��,A}!MTaM�h�MEN5E�*��<���hV���.���婤�蓒
��?�+��1m���N���h|*W�Vjl��ԝ��;�@�/$D�F��%��=��)�I[PR��!!��66�>��;�MB����o�Pw�4>^�ML�ء`E�����v��ˑ���x�n��Z��8��혤Z����m7�=_��p�׻��{��iۣS&��%0����Z��c��){�-:��D�@�a��^��	]!���3-�6!xO#��7�.8O�Wn�eVH��j+	A%e�~� �b;Y�J�
��a!
�GǕR�������#L�y��q�`���N�~�')�� <+����_7sd��Ɍ8��� ����Ӧ%� �復�zV`qf?n�M9&H��j\H�B��MUC�5bl���eծSS�v�UӃ�^�-��nωUx��k�N���^6�UT�T���u�
h��x��ǃ��.�>$�yV� �0�_�ʷ��̧}�4O���D9Q�va�>Ww>:Pр6���O�n#�hq�Q�>�׊��jV�@آQ�Ɂ6ѫ��b�����'(rNǯ����]:AP�Ol�ٚ��h��!Ѫ��:L�P.S�I:�O-Nt��-a#5��!��M@�N;#-��=��P�O���#�ӌ
_�ĸ���#�O�n�X���;GXnj55��8����~��U���^?w����B��w��	�л�� ����Q�Z�'n{ykG"�f�k��Ō]�R����vp<̂�=��=ᆛX��/�X~�L7Y�}e�c��ƈ"��
v�5K��ը*�q:ݒ_H5/�h�(�98,�����
`�ffIHjoy"E��<=O��s{�R��H���vff.\�����ꏖ��_�^���a���0\Z�R�7�"p��Ӄ��y��-���I&T���<}@Vs����n�[��c�C@�h���Dv�=q?[q@���PVn�p�,�V=�'x����x�۠������9���V�����9�'�Ϲ���Cm�ﾜ0gq !���[��kk?D��(@�·V�D���������_r;���%�"	�I�D�ftT푪��kh���5V���-�vz��R[ʏf�29 ���G�P-�=�'g�&������2�Dk�O62V�$o��3d��O���4�߮�h5��U��dz�;Ob��g�
0�F&�Gp�	�r��Be��"���m�
�67'���':�-��;�?�D;������5XOԶ=��Y�F�^�tE���������À����h����7�٠Ɏ���Ɇz����2�(m17����C�n���[.w&1�k�f�Mh�.X�f���1ݿ��eh�Ȇ1�jn{o�e_�Pff�����6*BK'y=�97�%pO��HV?�m���A�����S�bo��{��Y=���aݝ�"V�������E�EdJJ���JS'w�_{\�?�S��K�c@�YO�RG����N�"���2�+��%���������nO��*��0�Q8n#ë����}d����@��N�TI���߀՛�&]�d#�@�9:E\�J<�k��P�r���SV)l?�t�J�����i�`#��^g窜�d���s,1gϸ�����wn��(�Q	֑-�tq��B���`ny;	�����G�kif#�A�������|�v��Y<qόi��hW�d�����n9�����T�ҥ�����c?Rz�VJ��C��:�Z:*�8�>p�h������������:Z����Y�9/y�qt}N��#)\�I���sA��+C���M�/��1�8��ݜ:����8� ���KCh{��.	��mN�ڿ�ԓȫ�r �JK:R�g�&�E�J����jg��	����n��|<;�V�M�j��ng���@_H�huc�)�Ӷ�\���OZJL-{g'$ViS�u��s��[���(qH�~��a/�BQ�$a�m�2���?�T��4��~j�B*�N�w�� ��|��OB44�TW�W���FrwӀ�z�`��=�G���vT��{�m��X�Y�v ��������E���0��1�`\����ЕA�ٿ���Y�sw���ym���I;x�c9�&�(���z8�g�_��=�2��o�
mJ���P��/c�o�gM���?��������[j��ں�J�S��i�aRTp��$��(�d�U}�ͱ�i�M�٪$H� :M/��9YO��MOM!EV+��>W4э�늛:;)�.����^�����#��z�2�����i��}�����F՞f�2�6<|�I�FJ�E0D�]q]����o��Y/ʁ�EU�6�"GZ�F:�C�e���_����ڭ���2�+b0/��t@���E��'JF~�����(�>��5���a�Ձ����ۀ��r�!C�w�����Do>���B�Ѿ�v�T�S�]荷K���$��D{B��x��UGG�rSu=ozb��������3?��*�9qvؗ�Ϭ�� �`h-o����Y@����d�
w5�B#�;���PPgS�ө7��?�r�r{d�[��,��Yq�����9k�C_�#8�3
�裣���Y8\u�p�9B\��{���}SS�B��(S+��ՄAդ�Rn^�\^Q!`�����y�%`o��Ȁ��H��<_��z�j�!����R�� ��8EޫJK�}���{��v{�_������H�F-����l���5,`nn�d�G�/iU�_YS��f�n|	�G��rҿ�^T�'�z��4��U��L-rh/���R��ɉۣ5�5�9!@2�w9 �c�e�Σ[�b&ȹ����˝��3�s/��#��?f��������r���j��y�HL귒E�[0����e���K����e,T{F��H����Clz:�Y:�'}A�L��\���ѷ�>t�P'�������xyaGiE0=��97 �z>R��{�V����1v[��CDŅY�j�$��Y��q�`���2྘����	�k��@G�ch�ur��0a=P���%�a���o��<�r���60�uKb""��g2"������|ǃ���\�DK��N���7�@IU�1��A�r�w��E}Q����C�:�_��n{�v`��kJµv:O[3wmD1���u��F���s��d��g�?��t�]���$i�z��*0 A�<f��_u�Iw��+M*���3��*�KF}�ſK;�Gr:���h:'A祬�lH?/;�.W�.����c�nC��C����K#&�e�`e�2x�᭭$�����^����G� ��j�9�}D�,�M����P�"���"9@�T�O�Z�r2g	�����BET��ɮ����9�A����
��R֨��rҧ���-��o�im}IB�ݷa����S�d|N�U�d��F}�J���
��g��qڬ&��3= u� ���d�0Q[+��W!��2Ն����F����0eӂOrkf�ڱM����7*���xLi?$d�g8+���,��+���-��Q6�ͺ-�����I�ˏ݄ޗ��v�V�	.o������ݐ"`,Ks�$���Vƍc�` �́�c6Z��TbteU����5�޴��c���N�m۫<xv�qa	q�g�1܅���������2�uع0t�d��{9d��FI�p���t��0��u}7j�nS�<�M��������7�R�T���b7��ka�ग��ww�rV^Q�`�:�N�Œ܏�Ry��n:�y�+����FDཱྀ����x��R;��b�۵��e���ߢD%գ�;~~���0c��5,�f>�����I��p�����̇�`u:TN�BB�����P*͌���5��������mZ�8��V�d8�aC_s��`z�������eIvܰ���R�qF�Js���j�VHJ�+��jಉ{�5.΅��g�/T�0��H9��.����;��<�����04+"�T�l�+H���t��1�(E��t� M�
H����A��������K�<1yvޙ{��;3��)�C�%��<E�e#'�8���8aR�%��p�&��rF+:n ��u2�תk��z�<Y8G�zEEm׉�;1��(�9)��i���X����G���=E"�\��]�UK�'�l��.޴�7(��9�88XCB"��k�s�K��Y�i���<*Y.m��C�� �x"y0}���Z����Pob�{K��{J
���p���#t9�@b5g�Ͳ��7$��%��r�~���<�II1,�8 "F�#��ĭ�<O�hm�w����\Ά2쭞��sl	���A /�.����S-Ʊ�yĚp��o���x�F��FZ>�e#�(�N���D��@A�2^��%6�oLbk��W15�]@76��)�����ߛ`�}�8I�{waJEzv�KM\X��y8�PSC�|�����������"��{�ap�M!Rh{}��cK�*zyܯ`��`�6l�=��h����V���O��4T�KW��S[Uz�}0���Z�Ͷ��F��\����g���Ȉ��9O�S�V;���BMήG�Y͗
�b\�����B�l��)���.e���	�d�~0���W�+����?�c�]��f�>4�u".��l��/����D��Esө�c��BY{|�n� ~I���V��N�nQY��6M&&�����C�~��8��i��Z���Ы36�t7�tnY@5����m
<���F_4�w\�捖t zN� ԕ%���{x�ۦF������Fb�M�� �<�=�%v�KRH�v����$K0��P����|5: ����	�"Jn�}�ίB�Vo�%�D�FF4�͓&;��c��b�a���v�${�$�X�g��E$���� �Vz�������_�NQ�����ݜ�W&����eNY���Ձ��ӺD�C��($c(A���e���3*��Rw��W��;!��b��2-ҷa�4{�xX%�$����Z�Dj�f~����V���䎼�~��|�R�����+x꠼�J���%��CM��~|۲�5O���๞�����ɹ�8�7�w�V�6�9ρP��уM���cK*@b�\�޶i�FX���������e!h��G��g �а���΋�~����\�t�wYF?2]�n �Cw�� ������Nܡ�BAT��è��1i��k?��B�4�`[��W�S�VX��ş?�DϽ2޽��w�����%��|,2j���w�7A�4���S�.���i0q@�忴��ʋ3����n�������U~�y��rR�?�u�<��tK86�\́�� �ŠF�qG�/�q���Iڻ�Ѫ������b�pY
�i���,MH�����X�Ngv�::8�Ļ>�h#Z�c(`Svt�ԥ��͗rv �Y9����1�-:6�+�Ӝ�֢�Uz?����0ޟ��Y2�K/�;.�=&�.JJ�Q+�#���r��hW�:*\ĉP���nu|R��=��=�cc���o�'�J�?w!{o��H�YG`U���R����镏?�����;̨���g���z�6B�6t�3$��A��H���zA3 �9O�C�.��ď�њ����ƭ�p���}�^�w�ѣ��	7���~�Ue��BM�:�7q�8�M_P�C�(���z��_1�� �˾�����'G'wCf3ʤ�F:Kڒ�E�![�����әz����W��Jf�أl4ZAbS�4m��)�[����/~{m�,t1԰��DD,��� U��7lGߊI�Ӳ��~�	$�ݸ�b����B�L�q���É�)�$W<}�i�����	�������"�b�g,��Jk˝�A�"�BBaP���q��~�x�4ָl�������Uh��SK�N+�<�m�r�P:,���J��ԫ������O�o��DD�c��Z�g)ҍ�I��޾�I��g�n�l��r{zvFYY#D4��l�ф�k�%cÊ�S�XB���%�n��DKn/�I_9
�+Nc�i��79�v}�bB�ϲ�l��m��`x;hy����T(��~�$�c1��Wc���S<W7;&�s΁Mk�Ub�L}7NL0�	��(}\nQЅ=�LK�$ߌ����c���,�\Jܖꇬҿ/�EF}�q9���i[93[�~�mj:�{PԱ�d'7v�
O��1}�TDa���HQ��F3xz�kwg�����&�R5y���$%Y��D��(����R���y�E���뫿�.�hu���Yƈh���c4����Z�����߅�� Q�,�8�hП��� ,r�5~{�:!�-�����}�+��K﷋����GY��E�{�,�P�r�Z�µv�ŋ��ب�^|k�����!���{B�r�7~��a6 �}u��Wbj���2'��vᑟ���i#����ST�X�"b���~Sîo�tC��X�������jf}�lM��a�E_p4Ɇ���y��Ҵ?�N(Ei��U��B_Q�Oo��5�.0?��W236P9�C>�x���.�_�ca�Eu�67�i����Q�xz슼:�|�v�7�_��
�Ѷ�[�|��xVԞ;��^H�w���C���Ӿ6e1[m�0�g�s�P���M��4�1���`���ˁ{��l�ҋ	� �� vP^��	��aߠA��K��}���8�8�Gܹ$�^rcB��2�N�� f�u���%h>���EW�a�i׋4p����Y�G��^�Ǯf-�T��������}y=�,�*eVQҟ`ө���q�$���q�w����@�����Bm�
�l]����d�%n����s�COA�����8Q����x�=<�u�����\'��.�	�JI���z�$�t4�5Q�_p��!�=K�|���W=v�K�±� ��cg!�]�~��AA�����B���6�y�V���w8(�Z(��V6�额v��ފϵK���K�Y�|�1Rػ��ߎP��r��&��P��<����갈E��[�t�wD����I�;�jF���yc/Q��`+K+2�h��\
��.���r�:�`��Zb�X���ŚTib��xgB
`�v[VA+t����]������@��$*��ǆ� ��#��.��.��準}�M�!hEޒL�3"q[�v���e�G?�D��on4A��V2�(�qlY�c�(��H�L�,��]\�֬���i��¤z������4ɫ5T�&��wYD���:�z��O�W�l��>�P���W���w�S�I�NPV�����p�)tDu%+��!�}�F���l����9����:�C_�p���Z����z.��n�J+c��ӈ����K���y�h��
�'6�}g����@f��������=9�K�Iv'�$L��e������]�s��SB�y��v�E\�7�B��wJ�}b���E$�4"i鸳�O�r�������Ob�:P�����B��v:��K�	��@��7�=>�m(�&�a���6@E�r�E�c`��U��������E�ӯ��h�B�ÍEZIc��RwG�s�S�En���$]�tjrD�n��Ŷ����=cά U_tɌ���&@�b88  q���Y�F08���1�[ �x|����x�;�-qb���'���us�Sn����q܉u�n�!dkϰq�~��e@�hlh���Ǣ_�l�!:�㝇�����K�8%o�x
@�����}~nl�!��L���'
���5x�����|a{SY��2��gP���x	vdа�	w��#�IJ������ P�`	�-ЗM�|�����	�|�އ�a�e���u����c/V�b�ޙ)v=X����s�oEm�6���H��]���aUA�	��l@V�h��o�$�l�/���^_�����b�+�;��aE�oT�B��zI�<7N��йW���.��Ad��V�i���ǋ�	2mHY3��g�+Z������
�3�,�;��I�d��N�L�b��j{��
�y�ڤ�^w""6b�������;=�e짤Y����*gAڙ/���9��J�d�
�ׇ��7{b�ݺ��,m�1�Qo�8��3$��g}5?�H���WRc�G�ñ�i�{�(�-�[��������o�h�q�����[F)��H�[����|�p�������E]�^f8���+t���M���,9�H�[�0���twgĝH��-F�j{"�w��B������1��� '��I�c��(��;eq\��zn슈�d߾�~�;߃?�z�J�=I�'�I�[u����F�XП�9��\Bͩ���g�T�ywR:���\t�K|}����j�7���[i_�/ǿ9_^��~��(U�߳�,ӉKK�Gq0���b]�~�u����:��k�]9#��P��Y�������W��}T��y�:)K�rDq����܊�I�pɩ)C��/�6�N��a����5��m���}�����(K��ݑ1H�1�����1���(Ov��f�!{��N'zZZ�o�^��l��N~�f�:�%�V���B��VL�J.瞇Ǜ��vvq�g*��abd�	"�����������/0)c�����Nn� �8��muu���J��׆�U��h}��W~׍�.;�z)���\����\�f^��4�;{C����;�X�C��xx��g���k�՚[+��{�k�n�̺!V6�T`��n�f����;�\��.��Ǝ9��^֙�n�*��h���k�:��Yп`=g�Mu?��I2�d9,'�z���/���3H�����#�Ǚ��E%( 
�ru�s�%6v4OsZ�/g���۳5��s+���[�Lj�}�kS,��dh?���&Ox��;�I�����ۛ����[[z����AR&t�_ъ7ܰ�H����/�t��%f��l����Y �/`E��9�}�DO����
�s�4�W��g"+���;�j��>p��
6���ٕ()��~��m��{E̋��y˓����V=�է�O HF>t��k7VBkC����|��lt$: �����⢞5=�^o��3��s�Sw����hh�Q��`D�~����C%R�O�I��SzI����/�wϊ�UQ=�?��c'+�$1�U]=����,��ie��L�E�E6g�To���4�ܲN+��%g���f�x���jT��-!��ِ�	a��C@b�m]~��4d���؝���[�f�㑕�X����>���a�m�S�Z�f惆��U�"8/8��s�	m�<���j�}���W/��m*z�.���{t��H�-A%;vT>��JxR2��;`�귳	ņ�ev�~�	�q~_���oB����Q�3�x��c���'���*]���#��s��I=��e��\�H��z�t�D�{`��qq5!���ƛ��[[�7���}1�ЦT_qZ�d�![ ���!:�F:�M=
�r�D���ya��{����b>p֤dۑl��#�
�K.����=f��*˗"l��j��LG�:Q(�V4��^i�S��s���j�
 <��rH|�r�y�
S��9�)G7��[I�81.���\�r���'��tXa�23��c���dLA��s ��@����_������X��P��CF������b�B��)�az�J"���ޮ]#�{�����)�Jzazz�;ү���1����e6zU���b����i�&��ГD ��I���,	�.$�=�-���tR��q��{=qU,H?|�1buu��S#�T�;����R1L���g���]�Nv �Z��]���;3P�.]:�>1��nn��Y�Ei�fxlF�������glc���:2`����hii9mp����?.FŒ�O�f�LHg�L���Q��<�J@��T�\���V�(��q��������8�
Б'n-��e�@��<�ttTQ<�~un�� ��\��f�O��.;�0 �^��YR��[/����BE��@>(�����!?�ʙ�X���`2p���LN]��-��R��d{JiΥ%�j�T�eS��[Kg��<�cI����gYE�ͱ�Gy	J�(���c�r������g�q�P6X�)�֎���W�e�o��2���'���
�h!�t{ʷ[�����ji)�|��D_p��2RZQ�ޖ����K�����1��s�Ʊ�_<Y0^;�B��rF�Ui<�.h9ʶvׁ�O �z[��H�ue�������@!Ʊ
��������t�����LT���U(,�b�l�uZ� Ӳ��'��S��D���e�Y�by=T�ʆ}M��7L�P���^�D�d7y�CK�7�-tL�s������*�p'������;�&�=�_p���%&g�z�]��HG�Ի�"��O=����E7<�쌉 R8�<�xWZ�;�S1��Y6;o�L/���^���+�4<�|O��ʟ����-��N� �(9ߖp�0S��vH����5�z�`e&������_j��E]��s�<���/�Ѽ���o�<9!I;���k�n�$��	~��J�5�os����'��Yz����O(p����J)�BN��+����iy��4�O��x��OcO�r�lU��'��3)��f��q,O+_z��������Df�{��ŋ���s����\�k����]&gr� ���u�8\y�I��۝�/�
���lw-31��c^���Y�l�kg��L�D5p}@*����'�C�>*�;��;���n���x$z�d�\��ރ�F����迟�p!�w���n3��N�jN�-��q;��--�X������
O@5�O�;�-�T����_�� '��?�ݳ�Z/Dd󪫫���������uV�Aa�S����[��k8�x�F_����B�}���
w��P$�ܾO�La�����KYpt_!v��`J�2V}���S`�Ì9�|�n�dkk����:wGf�ckѫr������r�>��+De�r���yr���ι���oPmz��g��Rl?������(F&8�Rן<y���]�L�P�?����)��%<�n|{>����.V#�u)3��������wc���*���0[w��H\��r�v�7�P⎟�u�x龳�qϣ��3���ll�f�F����������P3���n<<�{�>��j�৷�{��F���\q�o[�ך���0�xD�s_F���dV[�py��p�YeIx~��}L.{�c�+@�
��{�(-�]�������_�گ����U!8�=H�6�,*}��G�¤�5��72u�0��E@QY���%��d����C��Y�ɟ�VL��G����u
d�l�ɂz��FNm<���o�wv�Cf}��Q+��`J�L��I���c��
�����Uo�d/�=�i�4�?��m�;�	��$�ہ� J|�}�����5=�&Q��{�>$ܿ�K�����aݢ�~zN��rp؜i����hw��`��W	uz��&�dJ�^�	����9y0w}�,�ujj[��B�� `�U�@Co�����R?}�յޥ!lV��ى�����N@�̎+����f�N�T�k�k ��ԇ��1��^�R���
�z+�ى��Y��~Tbr�n�e�&x[`��j��!ڌ!+:2:Ҳ�>:َ�l6 �)��th^^���/�%�ZVɡ2P��[{��܌��q����FƝ�(B}�˪ߚ�D�����K6N�m�S�,m)<�Kφ޴�c��G�jl�P`����� Ս�zH�'�����\���:��%!7�^�A��5){	G�ͮ:g54�DI�F�i��䮍�,�s����5\�����>4] ��5^%S��̂9�k�\�/�~~��R\PbmTI4FA'm�`-t��3���˛��V�_��Y�_v��*��d?On��b
p�����f�ڙ,�yъߏ��u΋�0~ZIួ�_��"�W��ɧ�Ɇ��%�����p�&��p)�N�k�\T� ��L�Y�O�h�k�0����`����:��:����$���jݳ1�N�X��~���Ώ��q���S���hu��)�)j�hE(�XF\xc�g��d����I���TUB�o^�d֎��γ���&�4��tB�����q��=�4�D���q��;&�AfL���]a�&���׌�ǥ�����c�y��b��/������'�>Ѥ��kA��T.��a��m���mk�D��޲�#7���6d"�=Y�����I��|H��)�U?��\]���@T~�诞�2l��	>	�7Hє7�>��<
��R2�ܵ{�>���#4��~�`<��eq��+ O�U�����z.�����K�f^5�8�#���0U��}�Hř�h����l����X�M�9)�Qm��;�B@X�2�� �(���ut��O�n�X�SVey�I��x�X����'+�޸�1�%��'ՏBtXW\4��B��Y��B�ж��n߿
4m���1<`����{�0�l���:�Rl������=�b-�;[���� 16��Â�.��=���'�25--l����D:z��~ �t�+{�*�R"I�3t�L ���yo�n�"WA��Lrb��Mw%ŵqS�Yk"J8T	�����TH�uqTYzل4|�V��R�ʷ���N��������;�I۳�j ���<�P��Oؤ�6�	4ɏ �`�E2w�9�M�09&�5$�f� �/�x���AcU0=�KֿD7��Y$�T�,��31fZ�z�����G��T��Y�2����ۇ�y.֘;�/%��+���V?������z��cGPt�vɪ�f���E��^Jn�%���(��0��'�R�}#�x���4��+.�Z�i*N�7����̰�� }Ķ~@�t$j8�uu��s��ot��b����j(tP�
�����v���Y(CM%������l�A<���3���I*0����Ke��~|�Ě6;eXFHX�%=��:��0^��u��|�77���:�;�w2y����R~�}�=�J����/��9�Ǆ�&�:�����熁 U�m:3-99z<�z���,��I�}�3�d��Ϳ�l�D�_Α
��>�I��{|V'=�1�cEsI!�����SLv�=�Ӝ[<<ڎvksKdU�:8x�Ib� �t#I.���v���,���F����\�q#'?l�t�F���e�܋Jl��ȑ�`��JG#4�̴�w�����չ(�F��o�d�bɊ�2�PUˏ՞5K�а�N�� ���h�}����;�d�����
c����G*D����C�ڂ�ΚD����.J��:�(�7If��ZeЈ񽖞�`�G���z���݀$/T���k5Y�h�]S.�k��׺S�A��2��BS�����&Zd{|�@mf�p�t�c�7��Β�Za�2Y]|�kG���#��[�����k�Z�BY��G�=�Y�B$����?��rK~�@�g���]�9!:?���><y"I{��{��o*��l(������9����Z��[U5��m��v����)l5��������#�D[�/{guly����T�r�!Ŕ8Ɂedu$d�֥=Uq]���;���'�����(�c �?�
*��Ř��,����`c0���g�h{����6�J7�ZX�,�Y����Z�`j����/�O�J�B	ސn��NlO�����_�G~9vz�TQi޲1�9?���J��:J�c ��Z��Zk��@����=���;8Buz�s���yk�u�=�5�����2���S�5����ǩ�3;ĸ}�>t�b�J�Q�F���.F̊ X���°� (n����{*�M:�5��G=�������}� ��9����(iQ D��"�-;mu�Cgo�RhV�ߓ�(�9�ü�D?���vNn�̱$*)��k��y�n����ٓC���I����_uP��� |c��W���f1�/�~�@�Oy�W=�tg�J�5���)��Ϻ�=9��J�0�-���	��&ܤ!
�7?'�
^������O�.���X����R��1�ɝ�Ԙ�r�p\_��Dׁ�]ļz����}�S4N ��C��3�T����iL<��Kɟ�53��+G�����}��3�A�����n�2~͍_��ؒ�	��ۓU>e�������t2 ��Ƶ-�9YGM�VV�\e��
I�~e�>�2�g��������tKg�f�R��=��w9������^'��_ʌc&�����pL����<p�A򏧕2hF᡾ӳ?hg�=�����P��F�������|�:��<)JT��QT:�Qgu���ֈd�հ'�O����9N am� ;]�����y]��l��&i�t��px�t���a����
5E����OW��q9�H
<�k��5+h��>�{4�o/��Q�2rR���H-��2��!�;S�
~��f��d�7���ﲲ�j�n�g�
�~�V��+@k�A�駲uX<��gB���c��y�¸ǻ�y��C˴����Đ<0w.��Z8E[o{����[eC����	�<FX��"��3�?��H���_t��/����5 ��ޢ_[V��7N9m��z��Q@� ˬ����� ]�M�����vT���{�RmD�ZZ���hG�9�b0nyp��&I���x-�$�R��{��;��?����7@M�{ɟ�#�i��"g�2Z���5�f��\�d�\��1�pNR���7��'�s)�$�<�5}���ĸ6M��:Ĳ���Ѭ?K��>�$�o�IZ�\��E.B�jw�~�2�w�A�s^��z>T�8�s�.4�RH�S)�f�s��1Vso�`��]�����Zo��[ u����"�b�Ny�M��xΜt(�����P.���
/���T�&,��T�&&Q�O��(�};��fW���NR8�*��~�U��T5�h�p�$Q:۞&�3��c�݊�\A�<#�\��ҋ�}Sܯu5y�m�~�O���I���X�������m��]fΤRCw\[�I��br޵�z�Rr�����L^�*��׍@���iF���^��A����;��r��E�XO	����)S�+��D�,�����f��=R��A�`Y�u��ʊ�cIa���Y>����V.�XTt�Uu4�@m���)�Άh�*���$���t�a��[ź���I7b�|��am745�\!��0�!1*�f؇M� M�1Ԅ(�e.��"p������̢$�n��t�.)��Ϲ������OZ����� 9����SU--m�,��6�j�2�'�������E6{�<bWR��$TB����3c�!���mf�|^-ࣤ�{�yN�8���P��ռ\��ڛl�4�Ɲ�P��c��#�r����#��t�/�u�X5u�8���_0�9��x�tB�)���$��<My�tzbׁm��z��1\��o��y=�/�7͠Hr�������mr�2��c^x��˄.����ܪ[r�:�jYd��
�=�Kj/\��4�|���/5h��Y#���$�� �aZ	"�S�f����a�kT�����ȣ�W�ːj����&��� �נ�4�v�u�_�O
�q�7^ⱆ
�����ퟝ�j�մo�BCE]qmZb����_��0���t���R��-�n��P��Xz�VE�_3{�Bﰊ���/+�kn���-K;
|D_��X?V����6w]��2d+I�t��9��YG�t0y�U1)�W�Z�LcW�l�+�a*d&=�����$�%�������Ը�C�~�T-�+� j-]�L�e���G�/�9e�~��B{���1��3��,��?U���"��@Uq��>ˉ�����V!��~�#x�\��(bk�Y��W;R�xdU7��7�w�7�����CЈ�a���o�1)�܄̺�h֑4�Ƿ�"��)�v����2U�� q��^�~�Z���8tih��
{g��0�����яJ~�&R�3�&��Y�PZ]�/[+x��i��&i
�U�Z��:N�X2��.^����5���,�T7T����&�Oׂ�´lf:�I�f���N%�8�b�@�}�\ŗ3�]�ת������Y\Uf�1�b�k�A2IU����u��K��@�n�Hڱ��)Y㏎�M_��B��"����z�Y;���;�9J$#��%����7�W���V>5=a�@��뮉I��Q�ba?���[����z�x=��{��
p�R�X�p<�=-`W���+�f��k%�ը��8����`& 7�K|6/�a�u��u&���{h�Q�A�C��O)rV�9{���g�5	�]�B����<������z��I�Kܕg ����|�O4~U���Q��9�����*%5U����Q��JD�}�M�ζ~�E�0YB�2�0�Y�"����U3�_��0wD��.���H<��C�7n����r޼�����]����[���b#;��8~ Ϗ���G	ʧ���x^��l�Y�t
P��vZ0R�I��u0P�3�q�I��+P��Е鳓��;e4�R�|��7�)y�n��)Bmi+�b�p�����M��+��b�hS��(E?�W�@�2H�3�f��69d�x��T�m)quw��=rcW(8f��=	��saw�9��!v�ӕ�>���U#!�p��t��t�\�;�H�A���?� �Oյ�~с������ /:V ���!��	�� �M�� ��/:�K����er�	q�o��<��k����ʕ�m�1-�M�;�0��X��)����c�S�$��NO��c�V����,�8^���;TYc`���?I�l%)QJ86J�id��킧��%�'	/	��ǭ�t�˟9�L�p�F�B_�G��lx\��\�ЬC#��$���m'��vr��g�2�؏Lk�i8�a�3D�;;J���AH���p}�d���ܢ!tx����!F�Sv�/�q	I���8B�Q��K�����1��ܾ3����79HИ�[׿(�IQ�a_Ӡ�(��*��B3e��_	gg$a�@ө��4ŕa76nȏ-֙A(\_�2Fǂ�W��?><�ڎ%|-H���4e`�)���������E(��zw�ʿ �ϣ������t:�X~O�zl����|��K�	y� ��ǎj���}�f�Ȫ��9����Wt��xx�z�>�����>	�c�Й��P�4ZH�D��$S�Ӕ�v�L�+��T� �l�; CHe�26f������jH�(�=X�b��~i	I�A5�g}^*��~��i2�De+���Z�:#�g�Z�v| ��w�*���mm�>��]U��
F�D��ȩFG�c�r.���L�v�H�Y��Ҵ�n�$A˅qy"o�5o$k���K�B�m��<}l7��+.����O1�Y����\W���d�ڕH9N?m����]Ԣ��o��� � 6���E�¢��S����9$��=+Fɟ�G����;?���ݱ�OZ@�ˤ��5E�����B����]+v�r��;s���=�37��!\zj�q�!V��Z���� QAxw�{�fv��k�<h�C*hXh_����~��ס'�w�J��ì�Wd[�?�� 1=(�7�g[dϢ�6�p�j�|���ܵM�#��抭�f��e��JKt�,�j������ ㎉�R������PݐFu<(	%����҉��!!���`^��^+_b��/ժ!c���Q8�٭�Ns��P`����X����?��HR�+~��(�����s���ruU�`F�q���of�D訰�hJ�i��'iә� vzVA�돾�e�ȡ[i��n.Ls�GZ�_�u.�eQ�}H�Y������#����~�bͦ{B�!$v���u���<���m��kSe����{hv{����M6'4&F
��_�]�bg.}(AR�����2V�g�Ũ��ۨ���T����4yQ�=��yE~&�[OOl���'._����'輒U���G�k�bI�	����ֿ]�7�Q�F�D��8_�+~hS��>j�n__�_B�x*���X��{��|��
W�G+բ1��䕭$pQ>=,漨m
0���6_e%cbsP�t�ix��	���Z�c.dޢVk�p�t;�����(�#*��Bw�f��+I��8� "-���L?J�O%n1;���O.e�㭓E�}kr3�	Ð养Z�E�]۵�E��!��u�Yl���*/pvd�|�����Uҡà���*S<�Be�Xۓ�@�+�zz\��?�6W�(NB������|�f~Dgd�6��9�-�Ф֬���2�b�;��tĹEl��O,���NI�8ZLH@��w��f�H�4��j(f	(pY,����
��e��b�U���>5��?
�a���o�jYK8:ݕa?�l����l;q���z��G<
8�<�JH����,��!�z��&��nvV/rX��r�i�(�.n��N��RT�^N^J7Q� q�����X����y�c��v�,�T�^rN�F3�J��j!��9(��Kk�k����,,(�G����׫��	��.Z��D���(pPp�(yܛ����h��:5v�;%����\�[J�Y�z��͞��F��>���K�e�+b[z�U��L�������[ぞ[+�78�	Xg
%��p޷i8O��UX'���_
$�+����ιbpS�e@�-v�y�Hq�>���tK/ը�-M�Rl)_��w�D��G���3���� �*DC�dX�i�5�}
�ߑ��ӻv���@�������d"I���x��p,-e+�}�%7�%��t���@�M��3B:����/�2��&[�M�����ݥ�k��H��<��b`��?�3����4ڝ�S�6��/���[�w�2Sr��������i�������oƋ���l����~�M�S�Qɗ�.��$���n�*����M �c��ڳj�2��R*�)3�~�+������yQ�_�з���H`�	���C���_pS�znSƘ����ף Ni��~ee�)>��5�����Lp7~�\S݅ϑ��	�c==2�(4�  ��e!q�UK]����BX��C���#�2q�τ6�1��ץ�y������eFr'��eĔQ.#�d�LtR:�!�t��jj���֯�F�ʻ�����&T�v�K�-A��C�Ƽ@]��V�-u����`3�c�އ}W�J���C|�3e`2��Tw��T�O�����-�>��,򔌝Q�IT���.�[�Y�^�4�=��@$��ɼsk�EV%LɎ�4f4E#�/"�;�왻��T��,���L���>h�H��";�"ՓX�-B�d5��Bůl{�SR���^��h�� |\�?�u�Dȶ�L<Լ��
�%6#�h��he�*��0�VA�DMK�Rh��?1�I~�c�d��a+� ����3�C���m���5]ro�ی����F6�ہ�7��J*7��մ�A�y+��Kd�;�UV��:[���Cv����[-���l��6Y���q@kq�;.�ٿm~�C��V2�TL{&�(�5�i_�CH�Q�`�znx����o}}���'�� ����R������q���Ld������:��r�Q0��L�(�á�#Z�T8�Ax��Z�fߴ���
�d��]��� ����~.>]A����-��7əx�?��8^K�C�	�^d?����ٓ�1Ɵ�>On��2]Wa�t7�v��XC7�%����m�p�Y������K
��B+[S�Xhp^T��v==j	,G5��K���Ȼ�7���)K��� <����;i��R�f��׃`�׵����BipK5���J��"�UW�xee�
�K��L��J�m��'7^C.��V6�������rAzo՗���3W�[����kP�p�-� �/ϧ���|�uE�!M\7���x��8��y?C�G�����7�"W�֢(R�@[�����s�Tt��O�3�o-�v�.����?���c��W��ixz	�j������ŖD�0�V��n���R���<��G��O+�8�>��?J�F�a}ZV���b3Y�g�e�uA��������.��@��X�_0x�������8�tZu���L`;o�f[���_�Z������7�s��lf�m�s
��u�ض�"�"�DF؊���z�kK������dy��0E��(������3NE���F-\�����!��@�K�u�C�k5�%cL8I�w��W[��:}��֕�]�>_�����&��o5S�j��\ƞ��}���*L�X�,���&����W�FFg/�≛��+ywH�v��)����syĖ}����x(�1`��c���m&
�E��5�<�6xgL�����8�'�2�7��kC�C��:�R�u�_C0�{$=��Y�3��T�`�9P��ĀGd���h�'�a�D(3J�.g���q�^rn�}l:��Аʽ[���%Z�#%*�!�~Ҋd_��b�?xT�y�-|���N��J����+e����f�c�#�(�tP>:�_+u�~U� �ԫJ+z7���<r�:�1��v<���1m�.x���'�	z�{@�������)q�ʘq�B<��M��J�H1��O9�"�i�=���^�L`��9��������_�	F�>'?����L�W�KЯR��T�w�ק3�KL����=��ոI���q7D/�߻�~�Oi*p7L{jJ��0�pTU�OMk��`�p�_��������C��H��@V���rm�08s���!��WP��-%HR\A_����h#�6��Y�UR�����#�+e���C_����bu��@��c��[(K���GШ��M-,w��7���G��z�o�N���N��(x�:�}$@�,�%��B��
�V��0n��uBG�#h����\��݈�����zV�z�Ks-�<�QGEr���Y����_�b����(����{�Z	���G�@�263�22]�1�R������d�Q����732N8����yq����E�<Y��SY�B9]Q�6�ua�(�!d+�n��c�W���~jr&8�T�y\���E5o6��0��D��nd��4�5���'@�D���Jp �|[��C媟΢4�8��fYV�H�z� ����X�~�Y���!���G�mO��Sx�U:Da���3�s^���U�a��i�qq�Τ��r��jL�Ī�$܎hT�v�J�g�pJ��J�f�ػ���I�АL�oϻ.h�d�p�r�	��5�j�u�Q��1���E�&���\��N��$W�[�E+���g�n�`�W\؟.X���c�Z7=������^��M�uJd�Bb��{��G[R�9Uڌ�a�����g�����S[b9V�=�$��#Ѧ���CѸۋ�w����T����_��gD80 �_NNm���VH]��q��u�E�޿�#�D����q�P"F���P�[���
ݶ���L����)Ӝ���7�n�J�@��Ѕhb+��wǒ�����A�0/���#��?��:q!�q��u9��o��yH���Z*z���'[arڎޢ���UA�s���hiI,3���/Nr�&-���V!�oM�տeR�ra������fz]���~��B�QJL���Lph��=9�P*���T���އ �ߦ���&��u��Xb#�0u@XلQn=@��kCUV�9��S��y)[������G��iS�6�9��`�a�َF�ov�g�����X��Δht /�i����W|{���ѓ��U��O�`�t�Q�@<|F!j��ڶ>�@Ql����I��O6���yN�
��V,F����b7-�6�Urlڡ��Ș�bl=����2���)�0�)�f`���B�?��)��A��Y�bܯ�W���ܜ�����/�E]�׹�Wu�Tʓl�{yr�.x�����_S�d9�q�	@������!U�lo�rriZ�d���N\��o��j�A
��Ӷ�+y�}���f��.�𤕦6��P���4mA���J���8�o15׷ߘQ{����g��+B����f�-D���TuU��J(��~G�cͪZ��/�Ñ��*�w�

ȷӽ�3#{݇��El) �ԩ��P�I��6�U8�Y��]�Ԭ��u�7O#&F��Κn��x��T��a��Lپ�
j�r3-$1�e`�O3F*\��xk��|1s�j�P����)����W�9k�U��n��)^P!��;�w5w�{�8����ܔ_��=�t�pkm�?��ub�O��^�WSYv���׺�_��l�,Y�ȩ�pK%�U��@���-�PXQޤg��Kv��v&B��b"��Db����ֿ3����ן��X+v]���R��uo����������TQѤ�o�I�Y���O���"z���\��bF�I��DǏ��B�ژ����"-�}�|rj�����uX��]�Ol�o�ҁ&(���\wj19'��M�~�ൗ����{s��'qW���Z4b8|�<J�9<���X ��E0��3>�'D�t�If=���(_��D˵�>*���$�����+)X�Dɓ>N��goN����%�M�t����Ì�i�������`#��pYb��;���D�n!sdij;V�����_u����Ct��7��2��F䳦�4z��K������Є��gXTW�><�L,hb C�ĂR�EQDA@�h 齏�"
QF@� �m�H Aa�(�0 ��9�P�������z�"ל}vY�^���>� �n"���'�U@�ʾZ:v�%?��y��RP��O�WP��֎8`8<����5/�Η�㖜��'�_�a:ߕ��x4��"ںOf����{t�ݬ���o8�_=%�m��a���{�R)�ڑ�F���g�:T��(���b&������M��~]/��HO)? �-eB�C�W_���*������9t��S`���s23q=#�r��������E����M�:�W���d�<_�5��Dj�n[
�����X{&���c{�������%��,�oη�ǁ��Q�&�������;I���I�\H�w���|-@J�I�^�e~�Ț���F�5_}mi-6�'�o5Rג9��ۈ��Gm<�J�����d��x���,�Ǔ�!���ڗ{L7�ن��ʸ����?Z���&�����?���촡-_�<K�(_D��DSO�.��#,�:��]�'X�]����r%��ȣf���88�v��B����qX��PVN9��&������쩆I�0�}R���>���ށ���U˾E��X��E�5lv����������M%��eiE�ͫ�qgG�߁���cv��2�އ_5d�tD	l����ui���g�Ԝ�-E���j�W�*K���`�����.���S�/L[J�XK�d��o��� �6k���b��_��}5����� O��{��ek�d0�mW������=�'^�l��A��F��eo�5Aphg�Xm�0�'*�!]˞[�R�bd�>�Y�-̊z�l@��`�����}���>��,�_ԏ����gfLp�>�%�ī,�̙z�j,�ZA�/n�z 'Q�<��_c��eJl�hRIե���)�0_~x���|���=tl��ޗ�G��� ���]�7EZa��N����}�-y��:`��:[}K�} M�@�N�"��	�f~žڠ�;P���6}�}�4���/����ν�Ik�*n�+q�����=�l��� ']��_\=Gݽ%��/ᨹ8��F��kL�E1��d��:(.�w��%�l�M�� �����]Ăj��d1��fy��l�p�K��2.:�������U�����_�����w� p0o�֧��(Q� Ȧ	�����ꖼت���b��~����N$b8�nT��$�B`����y���h{�I��]��?�� �����A����3Պ�pG}�:�p���GŃ.Hm�8�� 4�F��+	w�VD������oF��׌!�.4H��3��{�|i/�S�j!V��)�I'�5P8fʔ�a�t���n�d����~.��b�X(��_۞����KY�)�P.��{�h4?�^���d��
�N���ehz%�pt?�|�'�EA�;Tc���M>��Y1���"�/�&&ZР�gao���ԋ�Hi��EL�?���DYc�;�f'4�
@ɋe�ɺ}�)�H������5�t�������������g���b���;�<� WՃ���noP<A@i�'��pbq"�jwN����"�[��ͳ�a��%���������]���/׌�����J8�p����K��F�����G9��v~^%�R���+�*;��W��N�f\��,�n�!ע* �_S8z�'��y���`=p(�b���mY����:q�*�/�����:�">}A��˷ѧ^�u��MU٧��4���?�M�iz�K<�~:��]�?E�l�,�HE�.�3�����2UZ�;�}z�X�����Gf7�K�jX����ʲk��	�3ypFx�|-������D\r[Oe���vԄC�L�u{�Ꮏ<:����^I���{(�O�m��9�yth�O>6�	j�~��Y��np�}�9p�0M|^��X.����X��	��?��(�����`4E턬���.�+O�{ ��V�VkBU�Nm��k���3��gW$h�ݶٍ�耤k#�� ��ϛE��޹����g�oVs�����065�0�9Xv#��O��	k�}��9 5W�Y�M�����.[��w���h�\r)�p]F��O�M^ �tw�A"���v�×�0#�P��D�n�m`M� Iz���T���0h�����Ur�HQp6��7�\wo�<�TB#�O��q��U6�����,��znE�_([�G�L�;����ǯ��N����paW]�G��	$ɜ"��%�;��g3~ʓ���K���eb{�p�숄��yW������(H��N�����p���D��ǧ�׽%��_���p�ǃ���|V�P�~��k6�/ݓ����?�ޖosd�5��'zڏSv�	]�s���v�����*�P��ۈw�P/����vן�_�zۉ%�`"Ur��h���x��J�݅I�K�vd��qw6	%�H��B�n���E��˚���;TE@�S�D��M{t<��I�&�V�����F��
����u�����#�J�����A�a
�	���6��N���c���k��k^�X��m#¹kǳ�XڂMBW��{_��_C>Q~/���K�g-K���� ��� �&�r	�G��������fzP)K��;D���A��a�9ɪH�q��|F����O��r��3�,a��3�"i<ǵdP�ZN���Hwp��(+_���=�����ˑ�7�oSqr���dm�+X�T�v����� �+�={5@"0?�+U��ܕ�,~�qy�
�,y����>�0�܂ů ��'�AcQ$]��ߢ>?)e��ζ���uo��,���kk@�� �Zܾ�����$R�B���/Yso��;��D�BN{������2Q4g�/������~Y<B��kO����GQ������ϧ�g߰:��?ڊN���q���ώ5��;��9�+m��yK������L�ܼ���n�r����R�D{������C'/�n�X�;����;����;����;����;����;��B�9�6�R+��л\���^���R�pE��͉K�..����쩝�L-|A�U�v�ԓ�z�E�b�'�%v��7���^�˭���{���{5�ސ�CGVZ��7l������]�#���gҶI$\{�LHw#ZY�c��YI�Q!���5x�H*��n�L����ZH������˓�2�F����H�݉yVf�n\���Cs��"+��u�_c31����1��59g��_К�o[ۚ�E��_K�NL9�ipTCz;6���s�؊U����չ�9�>7��\;�ҳ��h��Qd����T��엀�t*�0�X�Ŝ��>H��A��-g�t��-��5#��5U��ji��ġ}����ڶ��~700�Ԩ=ňgcx)����4�>�0�9����1g�,�,��Ф��ϭE�@eW��n�ų́�w�	��~^�۝�~�`O/�R��k���w�㛨ў:h�����ō���bK������:m�(�AJ��F���Z'�/���G|=N�̍���^&؍��/=7��Ԍ��^�D�@��r3�h�|��G��|�>��a/7�� \5������2�ǱnV,i�	[���p�# �m2�4�B��o!�����	��k��ԟs����;rK�ml����er�#2c%�R���̹�x����&*c�G���a�Ka(ֺ+1����u�-�D���^��v�z�ў�6[�٩��Z�}2�VIav��E�;̍�A���I��w�Qsʼ:��b��.�� �^ݵ�3e��p�թD��;i7n�X�pw�d�o$�NZ�9c�!+pv�>6
�Cvp韮�������y	�I�#��H&����VWt2_:��1����F��3�a$�Y�Q7�C��2��2!v�LW|� ��t��v�;ג���l6k�R`Ppg&d���φ[�:��������S;�xǟ���j��[v���¹�Bn�V�Z�l�dH�GG�9�82��ue�w*C�2O��p�3��qj;����qP�ZN�O3{zR����-��+�z���n�[�F_e�AO'��|.E��M�!n�K�M:Ag9S���F�?am�1�rN�α�8hNJ�_|�]bE��{�n$�������#}ֿ<�=�>�(�����ư�W� ��eN�Bz�F[�#���t{@�����,.sl�+Q�[5|#`���Vy�"�-���=���������ߧ"�=:5� ZX�$"���9�'�{۾���4J����nΗ?~�reB���pe#��0 8(�}��a��֩�وY����~��'�2ݹ�ΰ���7����C���|�餬f�抿0o��&�ٙk���[=��\� �u`7X����k���_�y'�>N�3�v�x�XH�I�����e����GK�ʿy@/uo�����pj�������'�_)7~ҋ��M*�՞{�-ӱ���������ý�䴁�T��G����(�z�c}����LR�@\�j��TK��LS���/p����������-�:~�w�����I�y�h�A�N,q6]�E�V�]����xt�ˀ��m"�/0]�T���70��5��&]��Y�
�|��&N�.9��Ck�mk�����dT�⦾Zց��Dh�E�ȵ�6�RZB*�+�?:W�vs�q�a<Un<�����0;�/q72��κS�Y��t{��}k!�V�/�k�w�St��$f��6�<> �pE�3�3���h�����Ў����3���Cu�[�����F��7�Gb�{ҀF1O�tmT2RʉM���Y�:�����]����뻯�A-X��?-l�w�[�ͻ"T�$D�+��.^���� ���T�����
����3�`�a\Xf9�=�k���و�^��@�*�Aѿ�	?l4D�_��/A��Al�{��!���ީ������n��Og粙�44B��	�@�3n4���jh�$y�������bi�:vƝZ/f�yw#��{��*?#���PAN�ӟd���KH�2�~5��ݯ��OJB�� C@+m��+�3S_��C�j�)��T���{��9T�=l�s��zK�P��Y�kՋ�����c^`�)��W�����b�]5Yr�C�:1%�6,�Ӗ~*���DC��
D�Y�Hj�o�_��xd���!ڿZW���	�G~s��'��a��I��NP9�'�h{�q:�h09ikg!�Vm@�=_��R���ݛE1�$y�&L�nu�3�=�og3.��A7������}v��kx�	��RL���E�I陏�i�0�X O�� Yr¯��1�¹�%��1�P��.|�}f�)����vZ�~�|�Z����ִ�*v;O�6h�vw�dP��5
���t%:�|ZC_�����80����Z<Y�A��e�zB?x�iwGX�7 B�yS�M�{ib�5�7X�@��}PS�K��U}?��
sd��4-���N������Uv��̼߂\h���A����I爙��N�)���ߓ��+0s>O^�M<��"��9���0�;W���#��фi��9���|�B��"���hL>�2`�E� ��S�A#�ؖ-��J������l�U{�#q
u���ǟ;e�x��A�l֠~9l{=�Um�Q��?a����e�]�͙�S�J��NF��D�O��z.�n(��:X���|�Y�M���>Y>�;f&��Xg�+�K"����O{d�ٱ_C����9�0G�m�H�����0ˮc�'m\K"��H���Z��f�/���j-u��ؠX���F:*o���3�
|J
�*�O5~�H��r
	�=�?Q�[���9$H�Bb�هC&��Tv��Ǳ���T���ֹO��c
�4s����/�fm9��з�F ��k"Ǣh�N��(4N�.�㏯�� ٻ�Dd�)��'�Q^�>^�ItJ}�P�;�^:d����.���m�ԯ��n�+Y�4 �#k�}[a�%Gl�Q�v�q�£�oY�REhc��=�q!r�C�|��[�`��Q�.����q�6Ŏ����o�q�-�O�q�)�3�H(r6���Ab<.�A�_&��z��˅���t���&�jBk�ܴҌ�?/_�v3�1���Wo�tѮh�<Y�zKt[��츽�F�3G�T~�_r��2�F�!)W��Ls�������!eR��c��n���p�:.Fa�S�=�/�K�F� T��#_ـ儼��w3�:)����3�j��L����)	}��"4�m1�:<9ܨ��ѓ)�N����Frz-4�F����J���X���E�}oh92{�N�1(����T\}|�6���K,αj��m����E��FUJ]�hP�A�t�k��{|�\�GP>c]�6���J�F�R��q�@n������c�}�{S�Y��pr���0#@ [Ef�][Ψ���G2ػM-L.�~�S1�u���]^�q���hx���p�nޮ[?�ڰ"�]Z���"\e�Yy;�f��<m�Zv+.uB6<���:6��+cl��Wy�xg�JYde��}�I���x#1���O������#����rb�We��.�=�/�<����U������m ��+�+�\M�@��o'���zųo��Z��19v)�P4��N,{�P~��X�r���c��e��ϫ����c�B^��2�p�I_/����©M��Έw7���ƙ�柜9�w�t�jA�L�o�O�3rm9�M1�-�\��NO&�j��X��oOx�L�o:���e0��U�J��� ��c�����}����{��QVME׮��Z����j~��k�\P7��FUM>�U=���6�H9Bp2kcu�*'����6��ߪ'���|!���av��v`�3��zˉE�P���5���i�Roْ=�	�&��A������#��ڜ_\��a� �j���cg��	%��x&n'ì�'&�O]`b��Sī�]�(
�(6N�c���?c�ާ#�9f�~��k<c�b���2~�b%�����a x���oS�bsŻ�:�!�z7Qǧe�{S]S�u�\a$4�Ӫ䔑fw��=cO�ZU����E����6|���
ob,��Jy�*{1-��}\�ݗ���B0Ҫ|�K��u���/��N�G&�;F���m�/uϫ��� �p���5�;�{8L�,���N�*T5ɢ��C��VE�j
?�������p��t��ޯ��_s3@�a0gR�79s��q0���v��V?��ԏ_@�$U�w����X8��3+����}������$o�V����AN������}Op���j)�g��B��������A]Ǽ�;������)��p�xu��H�~���/�H�:W��N({���(���ۛ��N��Cۻ�N��o}�e1�	D�"}6�(hv�ޯ� \����&�?ͫޜW�ܦxE��N����Y~HF��s�֯���;a�+7��\��Y :C��+rW������I'[�����i#��k�g�E`�QM��
q&:�
4�-a���\%a��i+t"����u�	i��J�h�$l�q�y;ӮwZ�?ڱXе���h�,�U*�� k������0?h�%U��I�|!Q��RT�����3	2��T��ɌšMá-�o\��+z`�'���b�Z��X�0�a�O�ݨ�<mzc��Gne�;c�dF����%��
�,�ыQc緙��5��ˎ����SS�bw�5_���R���7w�)1������,^j|�撡4�i��kۊ�9��1x\�o3O �n�i]Y���	��</��99��ƺ�gbL��(ur&0'�?��#;�9�k7�Qp �A<�x�\��=`R��>���beE]����[�2��)1�>r���.��_�W�ɕJ�| =����ޏG��j�f&d᚞�`���CC�T������8�#��t�V2��T�xv�wt�xX�q�KUE'8`��ܛj����!G�i���&?a���{��i},fm�N����F3(�و�]D�:�Zd�>��{Ã�;�	+rf�_nv7��F�*Z8��Z?S�@GI\��xȃ���`��R�&U��������6�8���O9�����5��%!W'���9 "�����t�	��|*���@W1�ZX�f���en\	W!�����Sl>N��s �t[�����M��T޻;��/a�\O��Z.OȞD<��9��0��U�<9�XR8;h���cI���E2�do	�h���D�� �n3us�ޓN�Q�F��)�I��U�"�����a#�Q5<��
L���I̡�����&a	��2��#���@����p��dt�b��w:Gz���8oº=H�M:ꉸ=�+� Q��!1�5�C��n��\O�0��#��v
��Q��+B���]���4JOy����==O�'U�e �\`b�[Mǻ�O'QK���3���P ^=1�JcxL�ĊQp�?Gd�m�wy��nl<��,1U���Hi���&��eW�m@��<e�l��X�j+38�[zSAB^@(�f�z<�]���L-��\y�{���C����M�����޶�gW�Y�$t��]�J�u��o�C5pvƵ3	����!��YeGu~��
�jά�C�*[�;��@��n��8��*L�fv6�(�st�7��{�R�?\���BܖԜ�f�ޛ�:�.��]Y��5��I�3gRZ~��t��������R�k	�j�8n\��E�نǜkl9�<�8hS����|Y�$%5/p~�X=-�d�M���OjT<  ;�;�Ie���	{�um^� K�x��/2�ᕹ�Xc��ԣ�rbc�q�`�ź�K�*O�M��EI׌�%ݻ����C�bT�	���B�vQEHr�Z�(��J��W�Ai����JE�%r���Y�Q?���!�&�UX#�1 �GWd�ťJ�߫P�����<���v��s�\H�vr�N��Tz$�j�&�7���_l�jdÕz��$& ����ح��q���N�o4U�s�qa�Dx�J<v ������@qo��d��NpN*�}�@��ݨ��s� � �!�D<��f�3L&�0/�U��f+Ф2��*�Վ�P����P�������%)S��ݳ2�N��*��XdJӃ��4Ω��z|�%ȯ.�y�΄[�,�#FJ����v)ԗq��M��*���K���B�?r�b��aE�:��ϼ�4-�Ï��l��6��U�A�.*��4�;tŕ�k\��feKd	��?�R����u���w��L	솨��I�������*��:�� �0M��ÿ/hN�����P��D�B���1՝��x/ɪ~뎃�K�%��8Z�u�X1�&�4�D
�X�Ĺ�S��E�04ST�đi
���� �u!��IS���=)rB���2$p[�758�[�mT��1P�����fQ7�O�C����z0����;�ô��?�H����Z�cĽ �j!�(��8��jTUX3��qj�/mHID��Ӿ�?Y� 8K1��0��d�;� ��a�������;����{�^Y�܆�K����Iԓ;F0�w\mFRj��M����������{�Ԍت!�������
{!/<��,���Ow�}ε�����-�9�5�C�
�>�LK����:��퟼��'U�`y�n�HJu�9�l�nX���zѻ�[qOR��2{ȓhIz�hb�O{�#�{�*{�H��ڍ�l��i���F �S����QHX���l4��D�"b;��3���ح�>-�f��{p��ղ�Qgs#��	ĺّ@�|��[��s���P�h���ȡ8�����P<'Qmv@�+��2O�I�wJ�ЇK� }n�����Ӌb�Dj_ݰ|��x@)�^���j�h]���%$��?�L� �7@�g�����l��;������sM�$&�D������������.�<�N�b�K9�D@d��0��Q�Вs�Q0�Ks����t��t��HمF�
P���Cn=_Hf7������=��@u��)̻	��T�E����:�kR��{���{C�#��H����J�:1��f�������T��b�Ԝ:E� eD0��~�U�4�.v����_����x\0x��HA�x���g���Lħ�b�H���Hl�B�������{x`M�Ԣ]E�Q�X��&T�>X 	�?׵d�+��O�b��5Z`�.=�mW4i�Sh��%y/�_UZ�~4)?�~����")��c���1�`|CD%oS]S��W���n8Í+i����N����-��J�����k4VP��M�H���E��`�z#6l�],�ݔ�ک_�����Ǹ��7����f3 �.+qvY,�ǵ��
�b���Ķ���K���P���b'��j2�@-ľV��-���AF�:l�U#b���+O���z�j=r\5�a�c�|U���kP�ͧ9�O1!B�.RHw��Y�T���r��.($Vp�t`R�wp�l�'"��6�\r��]�/�4e��3�$;NW��8�k��E�hH��嫆,�*��X���bJ�)T���7�������3C�Č;>դ�a�#>-�~����/�������L�@r�LS�Ѥ3Z���-!E|�Wz]�g^��A�ɭ�k�ѓr|1XG��@����rE��L4���n�bQ�;�Da8�H�Dq`d�,?t#D�2�q���Gy˅��P�B"SU#��ъ-��B�
�'b�vK<����A�~'�Y�x���bLM�"�p���4�/0�����*]�^��M��:��WI��Y�����9�|�7n���v����PlZ�	�E�)�����J�خh�!�.����u��@�Ƨ.BU!�&߃�g�=�؀#�����h��뎪��>���*�L����*g#��w�[~G�!�q _�O�{���y��!�#���(��]t��0�Jޱ8����Dy4�� 9�u v�W�$����/�&�w��k���,���"Ƞ��P'~<��	�9X��H�}ha��yɱX��73:�����x=b� �mF�?�y}��F�
@-��#�_IoC������l��`c�����GAZ���[�J�69<�ħ�����	bM/����=�&�pT��(�ina��=L3ڌtU��nr���XЄ8`�[TCSD�x�i��C���zİR� �*��s�l?��EzH`��4v!�=^����|�-�(8��oi�[�>q9�13��ճ�*ԙ��fe�3���!�� ml�&�ˍ��V�Ux+%%�8r@r	�K.�/���v0D;c?Ym�?��b�O��]�-�)��P�T����=��u%��h<���\k���㊍N�̃n�<��M�r��O�:&s;}�g'�_�ܧ��*�2�
�7���'�!�A��m�/fԫ���$e9���X���}1w%�I���1�О���Ze1�ʉw5��?�\D�,��!���.V���W�x��'���m�=���8��ꨶpi$ztQy�2�b�u�j���	�������n H@���Ć�T����?�A&ʙ������YC���Ƌ��W�[�7Χ��Id�i��H��'����
�Jv�_�+�:_т��s�N�W߄���2���箻?ps;�f��˞�_?�iX�{]���
V_�> ���"�]1RBX��|+��h_���Q좦#�eT���#3�����Wa���{�K��
��Ox�����9M�R�@R�.ު$9�L��ؘ���8��1���RO��1�e{b�`T���DM������-�>B):v������.	��T�~��t����.bR����g:h_���M1����J^����oa=;���7e��U�	�A;I���l����������9�x���mΝOgC�h����/�@��i�t�]T'�3�Yp)�E�ʳ���T��=W��0[ݱ��g߸��W�u6��5�Q�xSG�����W~���s����ݎ��ݼ^[�D����e�L���6�مOo�wk\���հ �H�8PE:M%g���^�V�~��n;�ݬL�*C��n�TNb�wL�~]�ޘ��g.�?�E�D��l��XRD?3E���B+�(3���t�w��y�a�
�[����U�x�g�;����sg-d�����B��W[�
~+^���b��}�I�DYH�p����T�,��f���=�+^̈��ln+�rg���s��S���f�u7�&��PnqX%��\�H�_�	�j�[�u*��i��e����*i,���P�O�7��(r�a����AO���)9�&�'N8t�e�}%z.���HUU#����O���8M���7{�q�.d���?~Ζ�r��ju�wy�E�<�t{��Ā�h���9#�I���]��G�;M2J[����S����)�M������+	e6ӹ7�6�i���T����In���	cnߌ�g����z<K���
v{�y�2��5��~t��!�hF,t��vN���xk���}�� ����A4r��n�ޤ�ӗ�~|o?�w*�H�q=���&�hh&��Pf� f>eD_O#����Ԉ��}����ĉ��w�!������ښ��3Sّz�p�a�q�b�j&~5������-����ə��S��h��%��w��0�����0�
��������I	hD?����,玳�N�-�1>�����S�Nhq��ʏ<�-��77|�9"�AvIi[�Ą��6����"|W��z\ko���W�ig��p`�gN�Ee�JͰnL����[%�I��c���݀��2�v�����^RzN/`C�qF}tq���	1bV�]�ճ�2x�2�<��)8Uʢ��ȼ�l�IXe7��D���Y�b��8��;�V����kR���ӑM��|t��� ��ǹ'�<ث�����5zt�K�E��������;_R�-0�;�iD؉ن�Bu1��8��tiLb12D3�bR��q�dh��Z�-��w����ƺ�:���^1D��eK�J��4�j�i��qـ�B.�����A��Н\+�XJ��}tH����&�ﴜ��D�JM�4�Q�#�A�!�Ik_�������Z�ҟX�k��5#(~��V.�=q6��D�X�aR��7�l<.<s���jeg֗j�H]�a��a��S#e�m�����Giq�{��4�gΛ�|��ȧ�8�5�]6�O�H�aN��ե�F�iF����){<�o����'Z\���8<%��L%ݓ�'��G�)J�(ă�NSN���s�kxs����M��2�_�RǦ>O�̊�3G�JC�5^_������7~^��S|�A�����hj|8kب��N_��i�3x�>^�ӕ�<��W�y�2�a��cՀ>�~;u�ߎ�B11��85w�1%�k���z��-.����q��x�@.�7c�}��P�0�����\t�_J,���g������Φ���~���ZCӭ��3�[�$�f$��ˆm��S�2��
	G��g�he�uk�?�.oz�<e��V��Y�f�}�l����Q�r����Z�9�t�ԥC���:5j~/��Li��7��X14���N�U���8K�l�����a�D��^޶�ja�z����Ϩq�Z'�Q������x�0���,^�{��>W1.O�s�3a�;$z.�L{sB[�O�]����Jn_c��D��F��N�c���dn;�s��i �$�]�D��t�3?IMm�5����'�V���:�C�b��u��޳O:��f6��Zd��C��E�*UD����\e���/ic_��#��������W�w�::n�S86����U=�[�`��M����'nz=��;������Ѭɜ�U[Vt�;+�h8*�W���6C/�O�Y�ki��y�)5z��H:7zK@��~����sgL���)YO�<ҽ�
X�7m3҇x�t5b���g�H�r����x��'&AP��ӎ<����TƁ��%�[��v"xؕSy�uiI=%��/�IQ׭���7U��,]�v�_[&�N[�j����F�&�;��]&���}��T�͋�g�r%�^����mf5g���҅�6������p��(�������2z��_Y�45s�7�iތ7)����`)fܙUV�|v��=j�it��v\�C͏oj}_��v��.���Ok�{L�59k3ئ�ڣof&�x�g��y?�Ꜥ�^��qj��.ѣk%����]u�<�ˣ�݌wО�i��%r���܀���	]<�n��GT�~'�'C�}��௉�Y�NcA��p3���l�^�?�G��Tk��Ӗ����i}u�W_��}ȇ{�K/fS[�^Td�����.��gƤq�i)����6���O�ǔ�jA�v����x`��
�F����w��4�׫�L�Au��Z_�TI�[&��{r;����C
B����i�dٴ����CXu��)f!.;vX�n���u�W�a���T
%�A��0B�mmu��A�|R*L�+�흖g7B�QӔ�'v5	&V$�����ĸ���P|Jې��N�9���47ϭ��B�"82i�:z��q�Ln=1��9>pI�ً��A�ͰS1z������#���Ǜ8�P��>x�X�t��t�Ha�Lh� )���#S\ǈ��2�����^Q"�˞��1߷�޼�����	��}�.�Yn���%�^��d��FI9ھZf�ս?�oݟ��1%�(jk����w�sN��Z~�����HuM�!���X;}BB�Ւw�?LBѹ�xV"q���7�.R_&m]�	�z ��J�HC��f��g_�cB�=}�fH,�Y�;nS���`1Z����
��i��Qk�m������`�X|��c)�8RtM��M�D7����qW�6�ԫ��;����d�ѺO��cv�v*�!X�}�����>m���c|���zeǌ����C�Fx`�@��� �3��Rқ�L���O�T 7�e��@�H���j��,%��O���wN�􄑆�[J��ќ��8_�a�vwS[��r�� P�w��O�n$�G�|P90t8:�y�����׽ 8迪�Ć��!���;?��b�
i)���d�Z_����1�r�T�i�pvӴ���/?�@s�[�'󴴟f@Y��4�G���hJC�N� 8��Qn��jd~����0��gM���!�H�6�ޛ�]w�y��7'�#Q�J㾗~�U+cf�|5`�Dt��nN���0�� ��j������@h	܉>�2��{�ĝO���c�-���k�Pa���� 5w��B���9����ѓxG"����a�~�l����X5�Zp���>�$���'�b�w� �~�5��w�^�72N���r��,�L{g�� �Z��z�%�N;Ih+��M,��5��ZE27�B��͕I�hH/"��9���t}��b��РbJ�y�'�A�ɣ\эJ"em$�'��!+Ox�D�+�x#���m�zQ⸷���i�Lþ���<��~�0��U����P�*q�+M�o���*gAOM<mکA�Fm
�m
GZQ����}���#��=1u/B�x:�L���?��)I��CYA�Z��:�쾮����9.�Ȅ��x��U�iڊ�R	�|�$��:� ���O�6]xo�߸�Ï�|F�SYF}��w&�Į�7�N����XW?�&����-���w�}|�9!:5tLc�˭�4�3:�DY�X�OSs���d�z8�(����@�~Y��HiL2D�j΢%��b��΋�I[$<Ɠ����r f�o���M$����bD���Py�����C�r�x
���ף�� O�~/mJ���E�'����@;����-��jmN�į�B(aH���V�2ӵ�Z �:�a48���c+n���!�d�n���WD�_�E>�-K���S�-�:Ϛ��-�����	��(1��y�S����bP[sZ�}"�Cщ"��wL ��w(�`�0��o�~q�L1~e�z�����i�𴓎"��(n^��%�S'��_�<A����\�Ͻy��?Ag�ヱD�A9�^S�G�:Ju����RPұ=غ/�/L�s�����L��4�CM��� E��ɧ��������K�o���PDhHޠ�'��|��Rb�}�{,8�~s�wG~��g��Vd� �nRp".j�麙�ŷm�L��ks���������o�)_�t�f4Ppx��O�D�=]�f���K�H�1;�b
�y�|@b*����r�Y�w��\��������!)�Qu�PU��Cż��:�K���:k�?a᠂�
Q������m��[�^������oy%^��ﾚ�Šzg�h�_'�����b�-� �y9��,��o�[�͖H����l�·#-A�ߦ7i��9H� KE�hj|��?/�?H�]���x ����{��i�Sa̋��_!����J�R�߄��3�(�/�%�
dI�f��/1h�3���
'�^�b��1���L=��S�C�Z��L�-@]�F�o��݀S��8EmJ��r�nҳ����lZ��B���1y�cXM���A��qn�D6
O�CK���䥶A�]t�;������߇*m�"�lz���ܥ�/)��׋�r
DU�� _|{��?j�7P��+7Cf􀄅�HT�]����4��~�qM�|R���2
�����P�� �-�zu�3�a��х;�y���-z�M����QP}��Eڀ'�������$;G�d�_�X��A�߰V�f���U�Η������2�.P:
*�;�%��I�˨٥i��bZ��X�Vޠz_�r�K��6��1ZY,}�#�H����c��]w�3����	R���/5s���?�Ca���6�b���%^9~^.Jغ���-��K��1*C��r�'��?��d�|O�����G�K)�F�'t�S��ρ#-�ߜ�!{���9��ȇ��(n�)WE9�6d Q��"!�w���ŏ��!�Rɞ�~u��qv�¿�Wr~�^�?n��X�4����Mƙ0�D��Ma��죋���p&5w�Z>^X����.�

P�����Re�j,�;ӘX��`�1\M�l�p�ͥ1ʙ�q��czm��T,]���$z�F�tN�>�η����R�]_���/�1��fw�\xUzTN󕓩4�=��Si�2�>�L�E��  �$j�Z\\d�kpL�S)��5�G��&q��%*Ei*H�<xme��+���vI]����Ћ
��n�D!,���|���X�XX3�vo@s-�׉����s�7������C�D@�H�
[?�G�giP�Y�yq���Przs�������M��:N��2�`�b%p�_�`�1����P����^�.�uH?�����_͍n����Qvs�m����HeJm�<Ԓ���W��y&��*���XH5��x*s�:�v ��u/�� ���BA�f�ț��H>&���"�\�[��6C�4�_:�8�mn���"C�8�V�C鞎�AG����E�dSp�sl$j"�X7p����X�!�u�W4j0���SƋ�C�t�j/pHã/���'P���?~gR/���#(�τKǻY&{���9�C�(7��_W��-NB]f.�X���O�4�ƧF�,�	�#C�	�>���Ρ%5�6ɋ���.�_r��K�6W�6�8*�ӏ�[��c�&��UK�'��y�]H,�� zb��;��b�a}[�ԜG-p�z]��~fڜa7e;�C{q&���s=7�-7�]��ҷ�g\�
ϗ��hR |�0����#��6�A:�Љ��#f��YɊGޝi���>.YB*h�g&�vX���D�
7�3��+�q��)����y'$)�4�{�E����`L�Ʒ���26;����R[��� ��Y��C�ݣ����RB@��v-p��:{*�4���_����ct�K�-q;��Kw�UA�D���ʎ4}�?�� [9)(j�JI�	 !`�.��i4���MJ~
�/-�����e����;`�f}�@|�Jm/{� �]��Y�H?��7��q�  H���־���7�H�R�Q#��.�ɲ���2G�=�z�ͦԽ:�/�@?��\B�~�j[W�Tж�$�3dnKpϦ�RNH2��¥~�TS�q6�>9}g��;9c��浲{u��3�c��l��)�P�s�~>7�J�͜�-O�z����{���\.�&�kw2y�����/��*8�?��>���G��?l���t��G���6�D���N��~H�����<���oKCy�5�9ͶMu9j#&H��6�FU���Q;\���(^�>+�-������i?�B+Ruͧ�I���X�n/�e���\�k9U.�yin{]3��d����D<opl5<-<��/$K���'y
��-��_@|��vU+��-�<,t�v����{��454TO��+��։#�Ɯ ��'���5�C;����(�*�v
	U��_p�/^F�Թqk$��
e����q����/3 eD�9���f���d:vZ��m���;R���}�]^�9դ�^Ȥ�5Ri�r?{�#�jؘgj��X�ˁpT3{5��|z�H��qenZS/�9���$ˁz6M�pL��ܸ���nB�\����N5,q����V�][q�vu%8;{���%d����bi�����^�J����ڋ��~(4Խ�x)�2�J�quLm��v�)Ԉ��`��^>��
�w�;��m�d�t-8S&�~�n�Ƀ5��E�>"? �?���%je�Ԗ��:'�$dHW��Q�N��>�:�O���C_�xb8Y�n,�q/m_Jb4��>1����R��W�n�ժ�N�4���[�p��<_.|���_I1N�zҨ�����-�UW#���Dee;����\�s��`m�B�������yt��qm����6�
YөaW�N8⹌�nj<|�ʧ�M��T�.z���Aw�n٩S��Q����V�G�V0�n��»�����d���T�i{"�;��ߺ�t��b�͌#�i�Ƴ�ۺ̞�H�� Vn洞��R�K&����ǃ���MU
+ٛ�D܃�o� �K"�)�c��4e�<%��p�UUd�Z8b�:�1�%���<c�[#��������G���<c���ItB���E�*�u�����+'\ E��磞�V1���.q0����=x�ў�����og5�yױe����[�:�iI�9�$��)���(�ˍ��~�v�9dB*j��v\S��C�⪇+ﺪj��ƕmn,�$#G�y�� � 4.�m����0�sa�2RvPU�X�k����<�����:G?�p�����<=��<�k�<�87�������ҫ1�@Ч+���v{��ԧJ&�{�y-���[�[�׻^;��%�X��~�s���U������\k(^���O�+)Ó�����J	6�0�EՃ�I]/��o��z�	�4�v��u��~�#Ovq��?�y���j|�S%M�;Ŷ��9uD����1]BjjaV�sB��(y�!G����x�0{��j#�� {�m�O��nt*���B�˼S�5������p���L�WӦ	��"�r6��"4x�����������J=���)��T���Z(2aZP�ٙ�J�Ǟ�bHJY�T�^dO�=��;�w������>��|�����?�Ϲ3w�E����s~��$H?t���b����3p͠[�C|�R�n&����ϗrf����#����֤�Y�'k>�t[	E�i�;k����{o���z̶���LG�zx��3�`3mQP�g���(kFڟPQ��{�=l����E����uLav�����w��=E|�\���0>�V��]��� t�>�i|RQilŸu^��M��� 3��5���H����W�Z$]���#�{:����a�_��.�S�[��'�L��� � �ׅ���t��^7/�P6f��Q����|�Z�	�/-/zn�N�y6�a!���`�%���}N�
��]x0�ňP	���M˛���~����ԭ�bD��|�����/"�#>�[S��7�I7��v��l����l�^�d�?`���J��E��S�Лα#f��y{ 8(��	�_�,�]�B�F�۶B��c��+�ߌ�?����<h���z��
�u��}~�&�nI^���L�٣U���ߚ�����s��RS�I]���{'ނ�K���җ�i�+�A����z��Y�:��C�����	%��w�K��kv����h�0��	T0�K�\ҳ	 ]R���)���ۈ��P82���#\o��Ex�m��2��z��9SajT��_I��m�B��js{��б�[�?�����C@y>?hzlb��g�U8y=]�T�~��<��	���u��B$���\�J��,�gb-�y��0'o�j���O�$�Љ��~�u� X������'՘���|����'�г�b+�XhD�)�ʯ|QZ`�Y�� K딓�6S`���LJ�z4��Lw�8�i�XRC�yQ�Ά�l����K?���c+;#�$��y��A �b��P��0%%����������AI����ATsQR�&A���K�[���
 ��S�EW����l�ተ���:�Az����aM�b�����^Iv�У�t"��&}��X1��o\�Dd׽A~P������QK�xE��G q9�6!�+��V<~����&%�#��S��<�0���a��6�]i �`2��2P.��Y��j{�I%F���Byվ���]���͔8 H��lR@ki�y�y�!󋜚C-��V��t���>�e|VR�yh˹R�x���w#"���<��<�����v��7�$hӍTr>y�_R�t�?hn�iܫ
,�F��5�q�4�V�l�Ƣ.�U&+��Y-AZ�7��F:���6�_��c^1��u*J�x�z���V�<M��
�������!�S����Ψ���/!`\u.,9��`�h_����_�";�K�}D�|��E~XNe�ê&�������T�������a�N�-�P��v_R\N��ܟ���e���
R�r�DHG`&�oJ6u;tTt�=�&��+�Η�@��}μ �g|wV�3��5��x�����*P��¼���2�%)3VC_������+ѹ�AMKa���s���2t��7Yee-��f�և_�bL'~�SB���ڒW~�*�[�`i9�qL����ҍu�b@�;g�j���#��쮈1;(���-lc�8)������\�N�aj0�OJjKYH�\�B_UXL�Á��ϧw��r���N���r�=�(("�u��k(Dm��b�K��N�@m'*m]EY��TUk�\�?^ԕb�?��X�{�R���+�FX�K�Sk 3q]�?D���`��T.l'@Y�dc�q����<4���m]�=]�+�Ʋ��FV	+��\lx��3������l��$~��4�I��@�l����b^N~Ԇ��1,�z�W���1Y�hl�j�Y����E�:�V���y��?��	���-F�y�A�4�<޺3�ﳟ��W	�^5^��;��`�l`�Y�	���?������y��ZE�9c�)-<�f~�c\8]���$|SE$�\�>k��#���PU3����Q�n����������A�S��BcQVh��I~�3^�4��5b|Z�~ �\c! <�e���p���R�������C�O�~�9IM�0_*+��u\���������"�YյH�!u5Ξ6E�|�Fb����"Ҙ��{���%Q7��ձa��VBmL�ɔ��MCT�0U���:�2|m��' ��%1c� ˵+>/���ޛ�eU�1���vv�T8��A^��P:#`���N ^�R�*�$� ��?ő�]���/ރ«��g:�[�u���sm>8 6 �Vt�"��>|
\��&����l���m���� ���U�ٷ��Yl��2��P��J�٥�nE�*��ف���	xRb&�.�@З�/�
qs�cR��H�f��������V��F[f�.m��'�C�1�m}syq����d�*X�y}�n�=v(����ї�	*�+Ũo�,�G���
�U��Q|D>�_�{Q�x�1V�#�Gٰ[R[��]!�����<�o�y���&�y��K��o!tN�=3�W�,�]��G�������|�*�����,]�equ�����WvhK2�8��U������ma���9Kګ��g�m��̍����DWn�J��f���0)��\�S�mR�u�b٢���v��L.�,}�X�`��_T\;�:�`�X���%M@T�Z<^U���5�&~�\���@�F�*{��nK%Fv��7���1EڻO�KP��7QA������4�ڬ��u��>׌�L�BM;c�5��|Y��Ľ���S�F|!�"g���@ꥩP5��3�vn������ro�g��,L�,9�DD��l���>�}�i"��Ce��N���٪�}��VPJ3�A<ѭY���ߩ]�	�����F��l�oG��w�i4���x�*��`�!I�V2��Ï��i&�5�|�g1�t�5]��3v\=�#�c�����@��ύ�E��hV��sޭ̸�g�nWqWūY"3)m�qm}���*�0k[��lB���1��=]i�*)���|)�Fti���Y�����{s����H:�ژ���l���/�3�L�����ըx"�
�?c��V������_��psd�uy$%�׫�W!���)Lm��C�s$%ň��}�q��<z��y�^��(L1zl�r�ӕ�� ���ۏ=%U@�9����m�הּo:��$�Ի�����W��uд�����a�`Dy���,|��8����M��*��cIW�0��.D
��r��"��Ct]n�<ba��cq���8�1m�yܭ7�L<�C��2�d���(�@�ׅ]�In��f7r���V�+v<\�$H'��0�י�[|�_�/�z��78�#���=^�T��ű�aˈ�r���Oa
-\�1��S�=�7Mu�N]$t��M��n�K�]E���̂����C V�o-t-wFg��\ي���I&�c�m���=fl��A�|;���/��ʰx�̈́�+�G(zDZ����Ʈ�!��Kym���G�7��%�"J��lw�����^�,Z(�ME�	���c/]J��I�DX��:p6�p"^}�[��U����a?�����u�[*��.�+��L�/6��ի@q_C���N�`����=J�7�_r�j��j��̎�c�:�������Jj���N���"n���;�����v.F�K���FW|<��K�W���H�}��:���� V�����&����HXGRd��-���m�0_���HXF�)�f�M����kI1�J]��;�w���u��T,ў��n Ԓa*��! ��7��:Y�ԧ>s�-�u Z�+��n�*>nn����v��	 d�%��K�h��ߦ.�l�t��#g�I%���*C�э�f˖��4�y�6��iE�ϡ��w�^	cB��C�V��O�ˋEm�9��� �7��t�>����9�u�����A�Ins}g��������`�С�R�8�&p�҈p��qхhw[?t��io$-�I ��W�JxlB:~�>��oj��~��6� 2T����O}��++�6�����m籟21��U?�Բj a�^ځP�\"�Ah���&�_��*��u�\��f���=�79��b�W�T��֠�S\���_��]h_������b !��8��j�@�Yӷwƺ.qx���;@h�G�Z(X�NcTI�l{\2�@�4t1?��y}��y��@�Dn������N�I[�7�i���h�z���/GPO�cߜÉj��HSI1���,�^�
�ng�E[Q/�ڴ��ϻ]�[����'�Ae!�{������nQ����w��iIc��F6�gj�H%��Hsݐ��ב���> �2 ���!�:�FR�Z��2?����C�Ŗ��� �>�K�G"�G�$�;�����hg��lz�]�d�b�]�6a����c��KK㖋�Αˇ�E�j�[�c�!��߄����Z��ŲZ���FƳ���H�OױE�#F����b����}�_9G;Ń󇾚�Q��ߚ@�IY��mU �2����yhK+�!0�mv*c���e�����A�?���!����Nי-�_2���cCҀ�{w�����+�ed��FI_�B2}ض8�{Bj�)��.OVIB�=W�gO�5�A�L���o�vL��/D��n�c��t2��^Vk�E=I�n��nש(6um�h�/z���>B	2"�@�,Tpr�\c�#��ʰW���$zt*��Qנ�lfatO��7��&���G��gl��|���M����pb�h�Q N2-M^B[��T<��KP���B_?����y,�t@��s����+��	��P�<���j^0��#Bv���_!���ā˂��K�Ϡ{�a�M�Y!g��=�L�ʼ�3_����& �m�}#�6��,&@2��*˘?�����-��2b�Q�HghI � @^V�j���D@���ר�)���_�Z]mD p������ ��sϰ4��µ�����+�s��h�/pr�)zч��1RXɎ�p��KV��^+�"�;���ا0�ǆ�n�p� H��c]r1���i~�T6{�Ģ����☖u�j+#��[H�aç�OH��譢x�\d���Ø�|^����<M����u���s��r�}��~�[ƾ`�E�Cf������k3v�*�z�t�5������J|�#w��b��W�4���>�g�3���w6b���}P�Of�������mOqX]a�^�o	4�`�⤹/J#&���@F��:	Ҧ��Hv]{ꂲ�M�����0�s0�?�ȓ�nX�ex�>�E�j��Ȳ���ai��=���t��/�Q�A.~PY ��i��3�FK����j�a?��r6G�FE�lފ1�����'��n��>�Z�e�LVB��������Fg1\weɶ��RY�6�L=�6��ʖ�D<F��Ff=�  T��Ā�#�@����/z�z���T͏���^�V!g	��̋��d��~�"1�np�x�q2hH���ԩ�_��i�$F*��όD|NWx�<�Ѯ�(�L⃘��F��񣚄��64����r懗�W�
�:	����- ��<2�i��14��[��� ��~^�Mo ���@��O���1�_�|SaO���Q�����n�*HRؤHS��ѕ� �G�[(��]u�E?�컼���:�?z8����.H���הF�ɕ?ڷ%Z�]���d�`�N\&�`�&��ғD�Z�FP��ʵz�����W�t��!/یZJh˯��+cL	�+{-�]9Ni�������!�v�./��
D��T�����a��@h&�ۦ�`j`I��z���%�7f�&z�k�b)���}��| L�H��ň��-�Jl��x�LIf̧��'z*Ǐ�.z�����?1�C�o��>�5�3�4�E|Dq��{�Y�C*��d^����*�F��d�		�%#���\��J�Eñ	G�?R�g=]����%�����ư�L&���!1����spf̷��|�^�m���C���c�^2[F�VF"%{�9#��)'��9#��h���/���PE�vn@��t����_4+�W�sd�)���M���G�	-4�Z��í�;{��l8�щ΀������~ʄcZ�݃\f��c�ܠ�]� �lBtY�^�1���C{�{�2�3�.��j���jYۊ�+=��!�/A;GS*��*��Cdf��he27��yx���2�Z�6���k�G�g�Г��x��Ht:}+u��ؤ�/3��49+�Q��V�ѥ	�� tR1�0?{BF�|~��̮�w/-}_F:�6�����Fڏ�R�=�pD�7�����n��=&X�r��G���B.F�`Y}r��K�v0oy��fgg�FR�;?O��Z,���Z4����e��6��q'��-M�7,�H�?�+�
H����{1Y}�z�o(5�׉��~�XB�Z�j���y��x��2Ԁ��P>Kq]��_ rG���t��xp�_v���d�5t4p���M�[�(+�����]�F?m���6y-����	�R.}�˷����(��6��zKz�� 鮂�<Pu5+�=)�ȱ���X�O�/Ͻ��8؝��67�+�s�`h����ݎ����#�Y�@��3���zt�\Ͽ�3v��_��~��[��%���@U��<%�ީՖ�衡�X���H����	$-+&��1<Z�I1 $��s�m�M"y�L}�����R	7	�_��2���+�yy����	�
8C��h0��b�?� 擲�b(̗Z��
P�YEq�!ꀂ���������G���&������,���XVAb���t�c k���H�5}��c�!�>o��@��Bep���E:��@ɿ����S��>���Q�4 �H�z2蟕�;��V�!�ד߭����B��Ձ�r��ͪ��W�@�|N�y��Xt�#P�y�J��Ϊ����D��\�#4�|t����F_T?Ot��̅�k �ߕ�)���dI���'�V� X_T|���2.@��iڎEר�����a����EK�3 �!ତ4�+�uk�Ľe8���{��֙���#��V0d� d�]�����t${Z��:���^MEU�[�8un���Xs:�Ջ��*.�Ry�"c���}3�����?`Tb�K⟦�!�҅��x's�c�RoH��.jI��,��V����iԭVA�u��n(�=.2k�2�\�:T%<� ����|������q���]�Kn
5���|uR��������!�X�Jg߳��"[�󬚽|���]Z��p#�z�.���ֻ'fe������7~�#I?�*/�0l�$I�s�G*sZ�ж|�/�mz����w�Tۍ��3�@P�*�q���|���f�h�1�_��RCR���d�ze�~��f�̣��y]I9<a�zX�][�gq28�m���FP1��5��>�W\��O����o�߮'ޏ0_Z���e�m�I8=TV�9���|��X��O��=��s�삋'������6vL����w����f�]�Y�P���e�vS�'ob���+4��u7N���uZHɡ]�� ��0XX�Ǡ���,�ʙn5}K�;,��M'|�.ZD7���l>�K��+���45���Ռ�.EU-D��!���ϟ�Ħ������h��u�<km'~��W�g�_b�r(v�uZt��歺��D��!W!Ϲ��*��ے9�W��f���G�q�!��z,�~��~�k�_�o�v�2���*x�^�Un1��\A
<p�Au�O��&�1!��]��!)�̙�s8$1�Z���˗���E!��_A��ӧx:�?,q7R����g�Cٗ�!��5�����{aR�e֢!v ��>'�:窫p\}�6�Y�$�hP���L�/�Q���r�쁬(��i���(�e݀/{[ߧ���6��2-�9�.�@�8��l6t?��TM�.?��|�yb���بݜ�'��:�e+�i���o�O^���(�h�'dP����6?�Yup����l�%�v���<��ݚF�K�}C#����0L��)؊1�ְ��2�t�!��3���n[�Rt��P����x�U���(�-�����F�Žߩ��@�.�DbT�=���R[�(b ����G�g+�� rd�A�6bʿ��#��sd[Y��p����@��^(s�ݰ���';����ӕ7i���Z&]��e����c6�L�!L�7�c.yu|�K�_
�IpO8;H�&w�RR��]u���.i@l|{��^�l�Wb�ǝ �*Jxա�=S�> ��:-�Hd|�A�пX���,���S�n�u��A���uT�"u�(&z(q�?~nz�,��|�`�⠽eXU ����w�,�x�G7������c�`Q8����|���huQ���g��i�8��o��� Ф`�ԋc6[�����&�l>C�����&�\�ͼ<rIg��qK���u���c�=U�]W�θ�������X0.���Wn�t��ݜ��(���z�����c�K��:� �������}��^�q��W�q�$�+ƽ�֨�OkM��i5��F ���g8�޼}�0��9=пZ�Cj���;i��������)-����� �$~�H�)�-tBr+ Y��̟��3��1v�0��i#�Q8���[�7��F���o�V�cA#}�����e�6�.�4E�X�� ?��1�MwD����d�O�]�^[(�����[�+����Zb$�S���q*�˽=j�(A{P۹F�v��Xi�,�c��ҡ c�f�^��ÍP�W8�im$5���2��rԄ��rY�(���A�胚Ex0�=fC�����2��¢�*�@*SD��ǴjE�Z�`��W6pV�N֫�-��~@��,y����i�U��W�4�fg|���E��a7#A�6���3��ǚ�c�u�q(��sh�F ��x����j0���5�9��|�ҵF��o��@z5x7'�� ��߀K7���[8E���S��r�%�cV����UK��s�����/��޼��r{���`��i�s�(�n
OԖןb��-e,��^
Dmp�1��؄r�j��=Ke���r6̨�wXy�%����8�9cQ+M�� a��@�����!����� MB��0�3�n@�� �������\L4���O���	� `�L#j�oO�s������1�X�clP�
�~���j�� v�x�R����oe�{���YQ�{1��-� Ye��N�O�)�F`�O,?�~�����sg�².D� 3���Qmr4p5�!5��dX�Ӥָ�F��N��%b��;��jB�h�;Z_ؽ;J5@���];ʃ�iR�5��@W�X��Z��^��j��W�c�é"j�G��9 ��2Şog�.�J����l���0)�P�r- Q���X���XH櫿?���&��P�V�RV�4fz�>KY[Y�Pbݺ�"�Ŷ��"�|e�8��o��
x2��
~H�4�!3k��ӣ�Ig��c���.̽�-Z
Ar`k����OB��-Ɨ�����c��f�3~�̻���(�墱�k:Q������&
+.:�?���-C�CGD�7�1Q�7]�Ӿ`���m�h�$a���Z*�xr.�d��
�|r�O��̸�tb�������:w�[p~ ��|�	������B�n��R���F��?�,M�حE/���|�h�7��A�e��٭�_�Q�#6�{�+���D�}��l:&�_8M����� ��y�}enڃFY �liU�~q��򩧫O߈;��r������Kο�pC��kL_V���Ő�8�p�3�3a�gZ�g����4����y�:Y�U%�E�7]{�ia�5E�c��y�_Z��D��w�ȳ�@�|�^���Z�M���S^�h�ݥ�|%�����c{E�S�_�[^RC ��(�,h@j8�����5��X�g�' P���qʓ�˞���Q� ��Tw��\�N�%K���~�E�6��c� �.��{������j*�G&ت ج�����d���1S9ț+��9e*�9<�.�,�N�ݥ���+;o��(��e�|r�y�L&v=g�f顆��]�-K(ڂ�*S��SB����}?�1�
`�z���bI��R�!ȑ��8q�HX285�SC;KV8�%`�9���qdl����5���J��+`�M=ʳ��/������=�Fˏ�����%�<	�*2���x���[��b����O*:	�C����m�%�4![�;����-�0Xt��P�iE�4[
H����L�}�{,��~�!n�5(�җ���aO���Г����$�
�!;��U�\��e�N`���Z���'� ���:�,�!�zNw�_��<��>&X�:> �;�4�N��}>��~��Is_���/|t�1��{�<��W��p�*������vtk,t�x���]�c�f�;��y��1O��@�'��-�8���-c����*�oG��4���M
���>FЇ�� �K�h ��a��%���7r,BZ�K}~0 ��z�$0?��q�_ve�94Z��X����+�^�	���3rB��z��;n�V˼���'f�&�&�m�����3K�7�i6�ԝ����������h��,�LY�w��dA���N:Qg?�`2O$�H����M���A��N����0��:���g�P��V-��6��i�u�0�����T.�AǗbHf�{�a&��Џ5��kӋ_z�%: Ё�������}Q違1��˳���d�p&n���(�<3����B����gԯ��՘�Eۣ��O&z�M�4����f�p&c�dcy]�T0Vy��!@i�MF_�Ͱ!�2	*Y���+΃V>�F0����'�5��:Fa����5�7z|v��B0ܩ��7���6�X�=զ���F� `h��o�T�[�(�~m~�L�߳=��;`<�\%E���-@� U�(�O@C��~��S�?�`�B��??6R3��6 �;���$Ւ�߶u>*���W�k���S��ZD�c��:��"*�SUI5��)m���3O ��;��AR��װsz���1 �T���K�C=��9Mb�ƅ���|=�c�;��y�{5�<�~v�/�� ��O������@���n����3� 3�
D�o�}	�0p]@]o}c�1$��Έ	�򠁜gҕ�
���X�j�s�5�H��e�s�Y����`���r1:���m���:��������'p0Oa�ߕw+ ��_���C�#_amZ�6������쵹I��~��اiȶ�
 �\�*o��g�[w�Z�9�,���_XII�B��l�T$���JnLZ��rꡣ8R�d��:�[� ��a���Pf� ձ��_4�$�<`֬:�aC[,cqp?g��p�Ij��}�SC0��Q_����z�� �������>���N�n�/���?���%��W��/��|!VT!VH���½p�s�F W6�����x�/ڋ�����
_��Tg~��,�w�Mx$���3��<��Q�k������8i?$Kʱt^�`�;cM���1� ��P�bS����W�)`�l����1T� W�f]T�1���@�m��x�g�5����U�(T�g z(�/z����X�Z��B=e=ق�D�z����S/�2n�j3��YM �yβn�ڹ�C��t�(z��	ڝ_�mcX~��Ƽ��-�@ka������&���ԇbG�������6��X%i}G�q��D6+I�s��H|�z��H�ʃ
?�_
��	�1� �^�v'wn6Ⱥ�ȯ�����
�� ڳb�AI�Nz�/������?Agx���40�UI�d�z���Q�XzȨL��X�:����=�Ҩ� pe�t���� �{���`����<��4��:�[7�)�����9�XhcWYQ8L�l ~�K�������$u����6���A�o>�K�� j��7(X�*�7�cUy�pz$ik�~��h�U_��T����~B����{D2 ��+ޛj��= �lNwmv�J���9��Qu�Q��e�	�eDjw����w�-�;6�+�Yk�u�0"<�I�D>`����rF~M���C)u��,���]u���<��[
����R2�L�U_��j�i�~gbp�e|��Y�]�֝`6|K6��/��A�TT��y��,n��
���|� P�.)α����/��Oy��l��`#�`#cP��׏�5t#�`τ^��p�_4m���[^f�Μ�i�i{�wC�>����&&�u�gI��?�J#���nݸmn�%T�@��s������H����Ot{w���<�OO �������&H!�=�˸}e��g.f�æ{4�����>��(�B�D}�����[��9�P7d�X y���/���
+��~냖� ��I����A�e����]̝����0���s�[�3u��У�B_n�]_d����R�l��,D��A�1zQ�9�\\7��cqN�<�O�ap�o�����_�ǻ���g*.�,Ԉ;Ŋ�| �𾈑�^�P��)]��g������Z��6su2.����i���DocK
�(��}��.�� �����@���^+e�o{G^��WaVfC�e^��i
-L!Hhv2lp��r�@>+��(2�I����!����-�!ӡ�I˩��L�Za������h��\�}�sW),֪A��Ș��-<�bR���U�)v�G�hw=s�]��Wt�T������A�~��Tť5���%�Hk��-�<���D��p�
2#�C�l@�5�J}v�z\�@�íY���kP>�����W�����}�v��3z������	0�"�<�"���i&R���ޔ��[&5RAeZ����;�9u	7��9�GF�[�P>+>A�-��sR�5"�_���PuO®Wo[�+]��;e��J�%!ƭ����ҵ�4�����"_���H	�������*�OL����^��&��x�<o�1u�/��}6��9����Ow��52�?���[��jc\<g�c��T )VG�J�B��~i+�ֻ3��{z��3�,��� �(u�Y�-�����F�wN�K�l�Q�m���H��ڂ���
���`���B�+O�Z�y��M��5�(c�D&���5S�t��CX�ӵz�þ�L���\���Y�26�S+M���uܰn�m�'��Xt{�����7��V6���:�Ţ���neo�����,��/j���ک}���>c[�ݴ�}�mE7v��'V��E��߹��*]8s�yI���]8����LsFS`zN� ��mWĐ��4|u�u�J�;�����-r�I�����CF<Y�qqN:���`��Q&~�)��-�k��h؄���I���yv��aL��T#�wh��ja������fY��C�>�)�XL�u���{A���:SA��ݖ��敜�=�;o{¯d�ߒs�]�kF~>������Mm��L'�3����,�:^�ZvU�5���-����PE
F9�-��|H���i�]���.��A�$�*�ete_EEt[<D�Yi
#]��}�	���T��}|LS�V3�ON�O�e9)˂���3��=hv';G�}J�imΝ\�<8J��]�~7��Ott��ʉ`W���I���g��Ԛ3v���ݳ��=F����AyH�ͺJ���_�tPqw���[��x%FȌ��aWG����:��?|{���ǉKrI0�����?��Xfv��
ל�K����v��<&�9�c2�0��M�17��	q�5o��$ i����x(���V�X��TS�1�퀟-��y�鋖��^��PI4C_�]���S�����Y���I�ia�gn�5%R��{�Xf~>�	�g74�~LMy��ven����V��� S%_4���)O�j�r
�Wv3�H��c-�����Z~D�{x������N"�6��OM�`��l��I�e��">���I|�՜�}_�y����s�f�nc-iTQ�w�T��U@�2l7m~��U�SA��5l��=��7x̬���Ύ�	c��G_Alș����A,{������Э:���|�Q�K׹C�]	���X ������ph�J�= ����Y�'�7��`�A���L�>Sģaj�����d*()y��Y�X�ucn��|�־��9���K|���N��.���{��4!lm�')��K�r��4�.�j�oi�!/����}G��Z��IG�q�_�x�M�*�/�#@��R��M��ח8��_(_f鎛���#Տ��4ݰӁ�@�*<-�+9z&�N�D0�0[=���ЁCY��s�oMenb݀䜓.����Ǻ%Q�ĥM��$���H�:J@(a-��D�ʺ�� ����ݢp�z��dVs�bhO�{���x��r;����z��}n��Y��ݕ���霫��b:��k����&���8og�������~���z6d�?,!��t�� 5�*���*��X�=$�a��c��O?����)��W� Nz��|���[*�kf��ao]wAڟ����hW�w��4G��ץ����������Mi��x�4t��Ȫ��a�Ks)�����ebG'�:U�_�ퟗ�*_���n?��u1��Y����[s��=��d��e��GG
�뺃2ޒ>�l�M/WE�����q ��uͷbt�<񝉉2�^w�V٩��I�E����'��S��� �M�x���_v=<�EK�����_�O��P���_#�|�=}k���]C�7���ux�S��g����S�M�x8x>ms�%4��F���k*��Y4�}��H�AP�v��O��v��~F0�(��3�{e��7��m��f��wW��'ؑ�`�!Jn�gzI���2� �Ybcz��W�|A�х�4��=�����
cH�.�?X�n���!��ۻ���Y�tٺxж38W�C�R�uKhI����x��uKe����o+�z&�3��� �+HďI]��D^�PR��[�� oP���٦^�0I���<-�]��������-8�3�`��� g2��Ot���/�#�(����x�Ľ_F\�wFʳ\����Nl�1N�s%������V�"�r�n=V�{���{�Xw0��X��T�b*������|��EN�_�A�D�?녰|]Qz*>����'?���]�:G@����7y��6C�����a=4Cv��Tj�?k��y41�?;܋���m��<�ޱ��}zc�Q+g���{�Y������|�����B����W���a��@�Y#�_¢����0�r�dAh��i�����C��Hr$�~��DHJ��S����	qA�	�Y�8Wc��Q�,|��y٠Ox�7	�����:vnB��s73J��7��pZ2JM
ċ����3��*��NH�2?ϵwZ�³묓��!XE�7c��1���\{X��,�'QC���8&ޮk�;�z4 x.3fw�&vK��4����86�0�Yҥ�)�0�	������_��ڋa��ǟx�1&��G��	�\��0k���#nq������׵�ʵ�գS4��˗���g�'[7k��8�XF�B�7��G������i/�P�ƪ7zE�j�X�7�_ �d�[=�����&��J�^P�(k6'������ņv+A�OH�Z��C����i��<"g��R��v�SO�WRQ���&6�.t֞��I<5�O�X3<��h�-���Pǉ��4���;K�Ӻ��U�����cSk~e9�����H���AI�B�E��]$�VU��[���������Uż����y1�)=�m�����ݳm�j<��<5�2M�?<�� ���7�ߢFrϓ[����(�'�җ�q�ߦ �A�뺆jQ(pΈު*{8q;��H�^��$�:�q>���8v�sJL���
ZxW��?�[��H��@��f?���NB�T��+ƛdP�
 �d@�����{G��P�)؞�f�z�u��?_k��t��o��6x��P �v��,��ފԇC=�����)��RB�r��P��G�.��Kś吞��{è
��ph�v�f�O�\����@�*�g��c���`�4 ���]+�3pi\�#TW�[�w&_�� �5��H��؇x�=�H��;DiM%Ep��l�b��4�3u���w؍�j�سН~�]/:��:�t�ǒ&u�>Φ�NR��T���c{�\�?��	f>�D������jΚ����CB*��D��M����|Q|���.�'��'��ӤQ�m�)q�����G��l��'�UJΗ՜4�tu�h(^b{�����|�J�@��B�j����ZW�oZ �<J��O�z�<#����;����;
b�CI4�F@��t/O`��ˣ<]�Pah��r%�t�qA��Drz_0LP7.����u�ۺ����ӣl�@{ʚHmw�6m�����yS\��:��:3��v��b���}i�dѯ8��)7T�3�v�!y:j��"voZ�l>��^3�?�W��c�J�^$�D\[�{�ך��t���Ї��d��8m�ݳ�J�mn��1���%�����w|]y:EN��Hn�p�W�������4'��?rO��vCW��ݕ��E�8T���g����T�3����y5�?7�94��iݘ���L��*׮��x9x�ux��S�9��R��F��(����CD}
��2J(��*��,��Qq9�,���&�a��G�|*%N�+�P��s��;��EŗD��L�IW������"��o`�u��U��!p<�zn[
 ��
�~�I1�\*�?�f	��H�f-�`��ܞ\��i��T<>w����c~��hK�q(�Q�BS��_���5`��z�,��~�]`��%c�,M>��:lb�y�X!����V��@��r;�V3)� ��&����?�����ުM��� �5pRԡ �X|��B%�e6�]�d^�'9=�R7_ޜ��ѫ��y,�OY�\4]s*���] ���ksR:�k��e�b[v=7��)K�$)(؎,�;ׂ��+JA�P|wZcg/4b����T:?z��O;ֳ#̊N��S7{t�zrm��Ә1q��tu,a#��VPܑz���C>�zn��@���} Y��˛��f��R�J2�yֵzXc���7�
�c("�A��p������ƽ��<<4�LXq~5��j-� �g�)5�m��8���L��k�C��x5�K
�'�C� T�v�=c�^>�����=��`}=7�%�a-�#,��bR�epJ�%�^�-_K�����
'#�v�������_�Òk4Yб�t�ܒSCJ$!��u�mAA�������(��r/��k=EA,dWg+��Ȱ��8�wv��s��-�#�a��ypw��O�>}�74��$���5���j�!�Ҕ 7�'�����Z���w���l��t���������U�qQ97� O���(n���𶒢WP��{��"膔��9���8��5��y}~5�W�ihB%�����G4��@u�j�0���z�r_�lѫ+��ܗ"�����m�8�����<;^���E!~�f/���^�z5�:a�IA�����-\\�IH�X�{h�_���z�h����[a�PU!�|/�3[�̝��oN��27��c��qx}}����2�B�7%�ޞ؀�$�t,C����]��q��n�5Յ6�,��������F�2��ſ�^͢�`%�_�B�����),���L�S�~]N����(p�t�^l ��k�B�R]�9�Q�ڇ�kk�_����q��ރ���駰�D�ŏ�ɜ���C5����o@0�$����z�X�4����cn!��R�lrjj�R��E=�Sq�$g��\��5\�Ƴ���7$�~1I~'\k{#A�kA�?�z�9S���#{{��4��p�vYq�A�w�1dQ��oN~�����a���\�>K���+)�����F;�>ˏ�joX��A�T>F����ܙn����2sTP��)¥�7��x�Gd��'){{�qb5���DD+��s�g3ܩ�\�j4�����~�삷���VZV步����_��]�����Є�C�3�J:�ZXוb/�'�B�i��t�ae�]w��l,�? �԰��J���4�Hl����[?�%.P�uy��G����9�s����y��*�a��:��){{�I��{RF,]ȷ/`�Fս �oC7�B�{�X]�sR���m��nt���Q(.QI�*+��g�]�nW��_�kء����50�����B\����7@�:���U'��1/��Ć4U�p'	`'{��f�,
pw}�p"T��[W�Ռ�_��
e�u��dv��\�.,�q�R\��u�j
'��!�:�R�4Z�ȁd��xp�I���p�s��咏�[���^��C�+����Ce�U��/E5��۟�B%�q���i�_*Ƌ�`�2�������#�T��Ri8"g=�ק{��FjO]k���J�{�-�o
�YY�)Ӻ�M���!���uh	�Yw�w�R�
�%ǋ���z��0���$B�V�{��������P�I��
������3C#��(J4�L �~��E��S\l'��t5E���݃a���p��h.Lu����M����P�7�^uDI��؟�Ǩ�� ]��l�6��.,l*���<�R[��*Q��FC�����=�"��m�;�.�#x ���P� s�۫�~U/��d�sZ�@�9b������Ъ\Be!�/�E�j��@F�Y
bG�G U���6�Oſ�Z�z#�я�La��S���e5���Ԓ��!?x��g���-�1��9�dhC��9�G(˥[6WS�<<�PO�ԲC�P�_�Ws<�G���/������D$B	Ov
YK�Ȟ��eߗ�����IO��I�o)����!4c�:�|�{���������>���y�׹���w��[����������;A��$h�B4����tsB�߲�̧�gZ]�h��������<��d)���Mh����;� ��k�>�����L����oϛ�m@�Ʈ��À5 F ���Է���S�4oR��D�����s�����&3?_�~�<i�Zd�d����&�%�E�b�n���2iD޷x��. ���k��q���۷N��%��ѭ��ss̓�z��Ɓ��<��,�v����o�k��5�ZPj+�IZ�r%�����ٿ���n(<r���G0���B$����x�ld���4�r��%�����������Y-����m��M@#�m}}�g��G��bmu���Z(({������k0_�HCn���C�g�5�&�>qk�S�����vv�2��\wr����ٜ�2��uX^��]����U�����x�����j���	h	��__��?;�I2ˈ�ό虔h���A/�n�ĭ�'�mssA��,B��G����x�m��E� 3x'w��D�5��וLb���`��c�D��� �;
��p�ϟĽ�k�]s͗#@����{�qS�G>�~f�σ�"�3a��io؁R4n�3q�x��N ���O�{������iw��s���t�͟S�t������rD��ȱ錄�����Ԍ,�W?��Z2� 朏8>1��۬���r�_��>V�k�3d*�k�'��߶m�)7�e���%���#�Ǻ>Ǟ�y����I���'��tR���	ٔ��R3����B3v�Ԝ $Q�	NNW�У���[�-/-5S��U�6��)s������תƺ6h�Q"hɺ	�6����Fo�\����	�5�:Oh�04R��8⬉3)߷>�D��\��c��)0���W�-�>8�zY{���Ұ|=ߺ�����_��V�=�����Z��UHA2�q̀���(��3�v�'o���6�=�R�V�d����Fp�eGh�F0b����%j~ V�B9��{^�@�*��"�vj��K�G}V��Au�(m��G5.��}���/��!#��.Tj�P�EeJ
�KG�<ƯDd�G�]Cb\7 ֕�,JHX�K`����9ڈ|C{����ÐO�;Mc�'Ҷ����\��i+ȣ���q�Abx>-b�Ǘ�d�70#C�`��	Bs[�O�yxd$0�41����F�/�4���n-��]A�	��X�WD�,�� {<�9�FH��.��-d�<��H�i| �s܁&tS^�&���H��cQ�	�?(�	��RoT�</W�XJc�"���M�H��&��Pu�;����WA5��	��oej3P�E&�^��0{�[�U�N�K�'a��nGD� �% <I���?��_b��p2jl��^/��K����sZڑ;��I@_o����x1�h�ޞ��FO0Ϫ��--�o'�
�����'�+D�pqb�Т�..
4�
��MH�T0�V�^�K��?KK��*���lM��,�%�`b%�=���ڍZ5(7���m�О9��P�ƍv�#f!������g���N���%���l���p���FM��0��>� ����o�t`�y�߫{�>��*{��m��@��� `�U"�{D����-<��n���3�Zg�h��8��f��J7p���<�n��Jɛ7���-�@����_�M��-P���px�����#	�@�d��11-��G@��|��Ex5���@+Aˡ{i�0����(�8F̗����˜kk����2ww�\��	5Dہ���������%�f�`�� �jڠ��ۢ��F_tzz�2�a�:�C-Ƌ��O�>]�f7��?Uu�_.4��d��E�Z�SPY`�N�^��I��Y��
�����Wϭ�[]�Ե��!�D�S~��e��֕��&/��T�P7�U���t7�+�ra���P��4�5�8O�u��hnֽ&��\p��>��76���y3[��||����n9SN�����✮� �������s"���X
PZ�e�0�o >�3�^UWU���%ޑ��\V�)�6�t�UNx��QPd)=c����~��k#���}��p���o��_��<x7$+�$�m߇��x��Xҡ��ru�f���H�oB����˪�+A�=�ba������P��	�$���9W-> ?��2=�`4���>5�HEZ�������W�LY�+��j~�RX}z�b�X�F	��0-��L�d�HIPQ	:/�&w39�\���q��wL�@�hyʌ@Ӭ�V�I)u�ַ��(� �����U2��fܖ.yg[�7�8�̸Z�r`I��xUU^To�铓z6	��##��3wuL���a7���Р(4�G��Z3�J���b>����c�nqC�P/�Ƅ"3��*�b(��6X���D��ꅃ��JΊ��d^�e�U[�6�L�l$c�L�w��b���i�T���������xU����C�UU��Y8�%�[�x9+骫�+g������H
����x��*e2�`c] 7a��gh�n?'��]�>��ы �A]1r��s�#������ã�%c�e���L�]�\�k��	�A\_W�-� 9��`e�{6�,���ήO-;5$Ԝ�b��j���:}��3�?�6pE*��c�%hȤq��t@d�"}[��8���=�6�w���a%�s�������{^y�ME��G$IV�63���X�����]�Lrs��IB�≸���g�4�]�W9969`0/Y};؋���\i�%�QA
�����p�dL�ߧܼ�,���Y�Ò~��x^E}����������DW
#EO'�����<-���>1����w�I�j36X3Q)C�rӁ<]����1�}�v.U�L���J���DO��oo���
��(�W��"$f�	Wu�z�uH�1 /3�r��� �@[Q�l?�����I/�[ f�c�>�d�Z�����mb h-}�g�P��`�&�H��EZil�\�A$�hvY�3�<�t�b�}����A;�Ryv���ev�ç�����C���.�F�T�)�9%�=���N\��8��W��:C��Dw��tv����_��(�]v�V�
5.�p�+���r9V;�����:�} �OI���W!ݝ{o��f�����5���B�8��@�ي���遣|Y���J���qA,6�6j��틛��OA�$��j_p|$Ş�,���F����r����j�X�|��K|�S�,�6����w�M�����R��>�� ��w5��*!�!N���M=���l��|p����+���􆧾�E��,Y�@�����YBi]�3QI����~9�G2g�`�4ꕠt�@�KDu��\��������h��$2U\@��c���CH0��E��3�#"r�@j<�!3_Y��q{&��]��"�g���"�б�a�\���$)�	��e'����I��J��~{==ZU`N5+4t�K���_�� 9�Ԟd�~����	��"u]Z��& ���ڔ�j���I�$�1����EP�m��c�Յ�:��-; R�V��K^��t*gln��}��>�Xv�x�����_�b�AV���������N������u��fK��>��ur�EA���&葠(�q���ҋqzVm'��!i�i5A+��;8�N�W�g��ۯA!7���sx�O�>Z�:��Hۡy���q�_���u��{Ig ןIT�}H��qA�?b<E��P����U�~&������gh��9����2O�xA`t�i��=�t.�An2Uu�5�t���:�R==��} r���P��"�b����H'N��Z��4BF��̋]��K��C�f"(B(���%5�ײ����2l~�~�u�L����ϻ����-��B5�m@����������J��ttQ�8v�!aq��
��Р����s�)���t�v|�/�Iz�%�!��.a�W�gJ��:�t ����N�T�J�(XY�83��I�wM�[3���9<�xI��\�)�x@jv$�����=C�k!-ш]�6;�?�(�oh���\O��Q�ǎ��lsS��?��A%�Y�z�
 hј�Ls�)$!� ��M����mon��1^6��,�Bv�|����/���q�(������ɿ��+�I}Bx��۬uH .�D?,��#4Ck 6Ed��x�G�:/��$=&���cQ���jS�R��j��]�b� �.]���(@�뢥.]�[{�6S8&��˽n�p�#�h���R2org'�����G}�m��6Ӗ���*\����?3S�<�� �91����܅��j	��E"	���ym�����=bm��+����V�L�}�*����R

rmU<��\|p�Z����"ĺ��'�1�`�*Xҡ4��i���VQ,}-���fހE�c�c����iy@�L�oԈ���̂�D	�d�Ds����P�}!x#�+�?pn���~�\��ut/�h�ǾM��/"�� ���5�e�v��t!G�@���^B�+����.�@\a�����>�MԐ�qCC���OU&�3Yh1Ȍ�?1�sمf�p<�_�x���D��!Ŭ+q i��]�m�'W�鍘!�?�Ek6�MAT���~�8���~��A��ö��np(Aզ�?778VE��7����f�DCf�ۘ�i�2_�%c0q�R�Ǳ-�lN�<A�8A�0󢢢��� u�'���u�s�<Y��B⨈ӄ)�I[ZM�����>�숑K�d�=�,�;4_��F ?���L�9����[���=TG�6e+�@����WS�It6�����Az�\:�^��Q��Y�ʀ��>i;:Un���:r�у*+!�S����(�|HE����
�+�������������H/��pq���ez����(� fm.�������~U�̌��e��A�6c����$�}�{����r5��}���ˊ���t�>%W�����@p+7��Ƭp�밑Y�^��$�=Ӂ�)��� �3��{����v�b��FD�SdD���;/
y���<
7�����~H��T�B������T����{kOD t�~p�A����Ac;t�쟓{�뚗��I�Vk��E�*�"+�g{y��1uS%��Ǆ� �@�= ��Vh�>�����!��|�q�f�1i7,�t�.gi1�����3j�x����;�O�;=�{kޞe	���*y��M_}��(^���.�*7*�F���a�3H��q�(7P�5rD�/�n뾊Q�����ҭ���,]e��#8�ə����R�{F���V̯��׍@�!Z�_v�2p�=��0�+bϵ���P�V�P���S$���'а�Z�pe�g|�Mm>_�Y�!jHN��`2Y�/E��~�SRO^���>��
לMm�Z�I|a�-j������n�2��݃�Au/�؇	��j� v�Ji����QM�G���q�����F�T'TF�����w����}��xDO~ϫ?Ad|���jD]@�l���ܯ��,i�F�`�a(�-�F����G�gi�uKs�� g<s:�χz���M�T ʆBc����ڙV������2+��X�:������2�`���4���B̤�5������}[�=��M��$���4�(�(��Ie�D�HȆ`�nƹ��[6��b���Y�t䚂O}�?AAr�C9}���<r�N{�^�KT��4�d��u�&�Q+�'�n�+mq���TF>��N2l׬b$9��E�1�~W�l�ڭ%���^M~�:��	U�P�������@|�^�z�*��&���tv83M�+u֯�~F8��k
j�g��RV/���xس����ՖP���)M�g����_&u��u6}֢�@c��0P�c��d!1��>7K�<cJ�*��?=6�Ԃ�M��w�D1t~����".+{;1�@G"> Vn��&4���%�(�!�!�i��=�	{�a�6�y���p�J�肐��>��q���f�����X�+z�Lm�+��(�,���v��5��x('!���quT�8����r���?-�&�����#��&�GԞ\�-qJ�<h�9E}� |T�S��è3|����]¸�t	����h�~�j"�-v^I��F�¬CX=z,��^a��-ѣ��eNG�&��p�n�()�iԈ��#�Ñ>Y����3	��ۛ���IK�嗇2�!����'nfiΩ셌T�%�'�P��.>mo^c��ߎ,�����o����Ȭ������ ��};�[莪*ī]{�rI�u� �����}i��XH^$�*y���g����G��7ծ��j"ʞ�s;��zy��s�Trl�7MF��2�>*
�m�b%�u�T"���U�U��G�����3�� ��?f�]��*g��X+�,�*%���}^)���j�H�鞮�,�|6A��:fF�������|�KR߈cY�xDV\�?�P�A%�k�t$3c��2�އ:{�g;^�����⵷;-K9EC"�P��Q��-%��m
'<d�|G3'� -S�U���ڝ��Po�C���04f�'4�\��s���h�Q����Pm�a��`9�?.*���XW�N/�|(I�hKϵ()�B��Ó$�nT_��S^������Ae�����f���d^t�[��옝��ᜡA� v̬��������j�CL|'>%�ToiBz3U䏴����~�B�9'��ʝXy�p�B͎�O���}jQ��[�vLIQ�T�<�qz`��bZe1�h##�ݾT�L;��p5wrr�M�Ǜ��������$+'%ER_Ŧ>�՝-*������Jݵ+M�"dz!/�52��vWf���C{�C
�n��=�G~]�~��>�`W�T)HkU���o�5�wX�7��;�o!�#������u2����P����k��bRH'��f ��q�x��.���/�B�ն��WK�AnAi��/]�2�w��|�77G��
��'(�|�z�G��ج�k��76�s�{���l)��ɬ���hA�J��Nn#H�\�k����F�O\7��8d�L0s��$�*��� ��\f��^��?v¦2[-��(~�Og�)�tO������X�\�~�"�dD��&8����
P? ���b|�� ��=I֝V��y�l�v�3�鶷ہxq�BII_hp��JM�n��b%A����� ��I�x�	���2�K0�\�	�QTW�H�����\KUU�"V7n'mϭ�=7M���J�κ��e�QudTF��-�	%W��9�*(��֧�O���&1��f_	d��/���d��"��W���,;8��Û	�C�a	M�b3b�+8�$2�9��0�^��-W�
�	�s��t�́�\��#�^��Z
.�.Nc�An�A�L�g���,�n?�!�3�4��H���������Q�ǝ�D9�uKjk�]�M����+f0R���i�#��
H�SQ�~�uA��ghe�t
�3�j�s��g��Ig�l��S�:/T�tu��^sy#	5
3y�x�
q�ix3�ٌ�\IKgܹ�,��ʀ/(5n*���=����jo+���.
>S)l�`�)�WD��W����͜Ø�:C�W�#�M�W����rF�M�=}�ࡔ���-����[�Rf'�d%�$����M�F~[e
v���,~��#�y@NoU&7�J
�?Օ�>�9��䝮p;�y�k�I" R�ab��:E#C��}���q��
���!����ʻ�;��V��<h?ݍL���t8��:Dam jO�?��eekv�Q��å��yͲQ�}'�pJ�p����lX}������j쾿ˈ>:�h���"P�?t=Aj��p�[�]+3�k'�iWa��3<'��^̓?w�	����2 z4�K� 	#��sm��s�s�Z���nV=:�?L6�ܹK�3�l��'(����m�G^�$����C9NLЂ�]�yx����|��+�Ꙥ����{�٤O�:ҧ����U˻0�qf@n�$��OC���)�8(�O\`	��݂oF�V FI����P�㱁I����cGlA튔 (�b�E�p�8���Lyc��P�i[
yk_��$�@�ޤX�:����� �`�Z���J���.���:f&��?_��8�����W��g��b<=���Y�a_�djR�{㷪I4��abYC^�����;9�$£\�q*yok�6�r����_���ҷg]��5.���C���߃U�-�>�-m@��8�$:%��ep�!�*>3<�k_5�VB���C�J��|f��{⹫7$�v.�ٙ ���>��_~��#q���=H������,R����Y+��0�:c%%�kR���"��q&����R��V�ww]�5�K��,KD�LH�[切�e�{��&��`�ݣ5�G��|X
'P����Ư�{���@��Hd���C�R��l�HE��(�F����^��cs3��]�������E�]
Ww*�eS��r^�T������X��~��F(����>7�!���w�����Ak��O{���	����:jc9ˌ2��o��ǡU��O�9�c󺐡�k�	]���'�^^�3c��L}sL?����}v����ڙ�w��ׁ����B��<�����Vh�(�t#�	h�9�.���i���,mjT����������������e�0�����s�`^�6�u��k��.P&Z挄o(]��Xբ��h�:A��v#��v��k�h8�h��7a\y�g$!��Z~��6,R��3_N��;f;�XyGH%�
<����/��ݴ�)C�v��J3aJ�Lh�&�2�k}1SpvD�|>DJ߉X��P|���R��D��V�F���%��	ʨ�A�Y��{H::Yr��L�=��[/9�iv�ۛ0������yr���ӏd� ���K�
8: �(�.�D���z�#�J��@膦�v��}v�=9�����9�"-P�E%������<��V�$�;��ߍ -y@�.�d���XHXH������ѥ/cv����_�h_F,�B(I���Î�Z�I��,~�u�#'p�kХ�����$&�,G���cT��GB�3Kmnp�z:���<7���_]��&��'T(^M�/��k����#����u*�9�PE�����GI�F��`gCCA�ngZ� ���S?j�|��Q�K�.�Qv���g���[�g��Fu5_c걫�t""b�\Ei�:�t�킵�g9����ܐ�[t�8��}��U�>���RR�w�JO��9�x��.�EV��l�xR��m0�a��9ӵ��.z�N)@�w�cJ3���eR��<+l�:�Y�z�2�]�l)Л?�u8>��.#��g���zU3��>�MQ3r�nRi� I��W&�RgHڴf�J�� Z�������OW��Y�H
�����^���?U�	rz�U�Mq4�^M ���l>A����֛ޙv�����O��X-*���kY���Ŗ&uz��6�yA{�)wj�O3�k�!�ÍTң�>��� ����X��םi˰њ��K��Y'zJ��%� ~����o�ƛs�������r�~��t������ � �Ł���/(T\TB ��iuY�۳�����$1΁�_�F���B���L���JU�����	pHx�ZM�޽Xn�<���^��m��4�7i�/k°�� IR�1f�Y��0�?AE���������~���7fU��ɳ�-W9��7=�Q6���8	F�;��xڤ_L���&��`J��������ԓ�F_��Mv���F�S[�U��bi�T�E��0��h�A�aYQOd���@(���H+���Gg��2��5��uYY��,��˃ڒ�dj戴���b��\^�ܽN�����+?��Qk��F&ޓ�\�ذ}��"��an����(�:�O���������/xZC@"�t'V7�NqEE<-�E��O�hu^���ִ��%�z����:�]���󾑹ц�s�r�d��q7�w�DYAO��Y*~��͑l����D6D��5�՟q��M��y�p'�?�2$g�-.贅�(��=��Ͼ�z�	ݹn% 
D�g��]�����T��`�yR��R:��n�m}�_��@��!�B��Y�d��O�����L }�U%��i�)<�a�e��P��l�IՆ~��ڪH�cý�ӳ��js���H���uW���J�s�fSih�����d�'�'V�6�O:=�sѴ��Vn�gOH���S.]Q���ŵc"��\E2�!���P�D
1>T��J�	�7\QQ�tGyz�h�ط�x���IHx����D��<�8�Y;.���m��jY���o�[���Th�NF"��cSg��5� usS�ڛ:&th�cLG����$�-$ޅ��n)fҾ�1�}W�nx���u��oa3�����&Jؼ����qz���q���q��3kNNN�T���pu�ίB�>�'�$��t�zh�G���R�:�X� ����Zm�ԝI�ߢ��t�9�87����m-��CC�=Q��' �W�<c�8v�wC�-����C��]i=�!+{�E���G��PgC"���Y9k����ኃ����[1��Wĺw�����5`���Au+�����@o��UU�ɛ�roS]gZ3��(�p%:'^(yCG2;A�kT�W]���1���v��g"�ZZ��M��4G���u���O����gĭ��Bѥ�{�p����|T닢�4�'����i6�a:El�N6Vإ�~4�/b�\��}*(��朚��r�'���^�}T:;m���u�Y'�dF���Շ�A�K�k�%1zz���:����B�H�6	j�.u�8�g�/B6���<�_�	Ci�]�	yVp5y	1��$_V6Ԫ����.#-�{�r����p����b��*�7޳�)f��[������.Ǫ�t ����vA�Y=0y/OZ��YR�/q�M�u��;�ݧ�ٴ�#=c� �
(�Z�d*w���"�6}��Ɔ8���y�V���B�f]��S�jlj7J��!�c��kލ�b-B1=��(��@�t��p���n�R�´�9)Պ�����K�V������!���̀5ǰ�m�i�g7D\"���L���{��B�-����[^�����ٕ%B.�xS	�fݚg�;/K��K��6��&ZZ��A�2����&I��c�6ixkP��z��MW��2<D�E����r?���e2gj���� sQ��`J?��	�������==��G�a�'�d�1
����g�	���XHz���,�6��!LK��{��=&��3�{g~]��n���ր��޹��_��"w���hWE\��V����o�:�Zh������l8|��@
�J��P�	$�S����p�TTe.�.s�34;�Q}����-%"�����K���XB���fF���V�a5���r�lN}]4�R��5��gE�!�'�%C/͌:&g��_��x�{B�DE��5<eWh�$�-�6%��u'��V�E˝�i�ˎ_���W�j�3]K0s����D-o{��'�bz�>�N�@j\��ZB&J'��D���g�G�~���FY8j�<�)ФT�`+j�R��"ٝ9�����Ǧ=��[I6{3��;������I�l���Xj9ȝ s���ތf4�T>���?���c��I��^x�|��q:�
���� (	�W&l@3������h�,���mE��Le��K<�!?wN JL�@����t�Zg+���'p �*4c�<��-c>��O��"�[<�9��%`��h��Vn4�0Q=A�Y2����$�-_W:X���յ�{\4K���/֨.�M9$�g�G�gK�a��I���<4j{�m���a&�l�����C���p���~]q����|;i��ى&ݹ�\�i��M#�x�����~t*~<aI�B�s��5K��A���o<�%LL��%�����W�4�wD����E5��)Y�i�j��������vHl�>f��=��b\G�<�Q�e`�Emy�r{{��@妫W��G�G���"�@G�:��h�Y�"�&F�Cw�fI˥�վ��c�؃�
�;���Ƥ��M�����u�%�nyU�YA'X¦_R=�Q�E˩[5��g�b��5[�[�F?�h���=�X6�y7SR�;���I"�M����7�Ӎ����M'�xjgO,r.��s_�[cS�z݊�c�������E>V_��X����`Ե"w��c@=�loV���Pxv�خ�Ţ��-�n���	���^V���/�䓿ہ}�󳵍XD��T��ms��2�n���
���✖�If��uta��^f����`��?�^xTq����y2ZT�ΰ@��qѕ^����/�E��]�g�,�3�Y�vCٮ�Y���t�=�y�Y�qt�Iٯ�g'��&��9o����l��_T��)V�RhJ��4���n���H�L-�G)27s�ǳ:I��Y��I5?�YR�X�F��\v���;�S�m���k˽�����;9�C���7i�]���8歕)�w
	����]u�V5z��`���	BB��}j��Rô��+f�~@j���a�0�!�N�g�4Zv̤
�B1]���$,���f�����e����ە��XD@��]?�e����綪H���3x���q�/�.��)_m����͎-��yx���,�(��1s�Ǎ:+�C���K�O�Z�W$�F�*/�y�.�b�)Ø�2��f����Sa:����F?���q�G~��D��9>�t�M4�v���{���#r�	�U똩�c�ʫht�g�u1�x/����es�h4��L�?T�{tnt���v��W�%Q,��vo�N/Ifv���{f��;L��fVE���G�/��#�.����"�[b��'Zj��?R�\��_�c���U�* yKmj�|^h���L���U��I�&P��̊�}�7z!)i����Ì(���s�Z�z���7��uUڽ�o�3+ҿ�&�o��j�|×��b����V�u��#�������&D��nX���(����_�����v��jm/����LN�n�m[p�bnqzǏca�! ޅ鑹��%���������h�5��E�������$�Zw�Cَ�/�uh�qU����w�2�p�Xտ�����k�Ӳ>���3ή�t��IО����W�wwcS�,ރa`��dㅫ�j8������[˅�鞆0�R2r���Jע�x� ���x���s�+|�����a
�M��/�.z�ݢr�G�
:ť_Z��jǡ�eǼD���%k�WR�XL��f���)��e?��v�aXN�mM����-4'gM�L.���f���m�4"x�z������
�g<���vy.��E&v���{�X�o�"�
���0�SJ�]f�:3�8�[��%�6k&�9�Qa�|��kc�VK%�� M�_�0�y-7��CW�Y��)�M��w�����#*X)1���x(t�dЈlʉ�~��]���)y���Һ�3���wʷA���v��=g��[A���abڌL�F-k:��-~�Vqyy�9V05�Z>�:l�oG��Ȯ�f��h�O��=�n��S��R\���?e�;n�&>K���v��(�`IE���_���i�=��'*j��9��d�p�
��Y��.�ԯ��+�Soe�)�S����.A�>�:�p�Z�����5웳�ޡ"���έ�'-��蕷�rI U�O�{�*�������e�������+����\�v5Z[Ӟ=�My+�E�se����4ߵ$�?eEభ�1��
KI6��;C�睎��YF�=ȜBjZ�� ���~��
 �Ȫ��#̱�/�E��r8k��`G$Ѵ^(���:���TI0���F$�pa��b��]&GDd�$�x�����<�OMnw���{�^���z�sjΟ58y39�>�!22s����W`�+��b)��v?����X�a������e�������|�zVs��A���!�s�o��v\L�g�	������2 �,ƃ�l���š�����;��	����t���۞c��7Y� 'v��ΕK�R�7Qҷ�w��Z�I�<O�mɰT�M={WW��Ee��a�[�K_��b�>��y��DAH�<e��y�:�&=#��K�2��OJ��s>M�ϙ�.�x���9��P���s�#�; q�1,����KP���㷦إ�,�Ym� ��+ ����M`*6}N����԰{N�[2��;¹jtQ�f�-����}�B�[2F��V�h���2At���gl��;׍~m�Yu�+�2�	���K!W`H�[_6��EVk�Yb!���D������g��;�[��.����q9�n���(�H����B��A^�����I��=l/�D��^��h�cQM(�_ZcbQ�;���CٌOm׻�5N�'J�lm#��]�B��f	������4�`"@�#��o��8j����}�x������Y�W����,y���|�66��J{h��Y$���$�����5�� i���G�e�J�}�l�uk�4W̻�~����O�.�	�n��Aײ���F5[�z~�wo���+"8,t��e�7�_��)������}4�1�ކ�F�A<pP�,.?G�ï��?�8$z0��,u|{�|¾m�OR�^�pFb��(�G���<LM�.������L@� ��?^|d]����n�Կ�����J��1�(��B�o���QN��f����e��T���h�ҳ��E�]�0FP��Da��i	V-J��u�»�k��P�ɛcyN�Yx<Sb2�K@Y�M:�w�n�"!sse?z���l��L�0#�'��n`�� ��G�&����<�������߶&���4�h�<�̊�m��20T95��i��?OH�	�'������}C� ��h�'�s-(��p9(��gM�_@��30N2��͗F?�65GȮ�,��r��3Nb�(�V��7Zs���*�Q�U�F���ICޛs�����c*E�d�$iD�f�A��߭k��N`Ys�X��
�r(`�H)�F��Z�Z������X^^ŝ�&W�sa]Ե�p��T`�I��f�+��v6/��aR���O;bG�%�h�����`K��X��d���h?u�|���4�"�u��+yC�س,��Mx��o̝�}�Ǖ����&�0�)�$���^�ɳv�u�K���.M�D���5}�������gM���[+$��v[/���"�I��h��w]�}g���N]�w2$��@�Zu��P.:�wf3��b}@������D1	���k(QS��s{uOx���p��Դ>{�ë�n\.�����#�"3�#,Z|�i@���x`m�LJ�M�B����kتӳs���m��0X�A��l@0�aD�Į�0�~��0�[��7����Á�2S�i�&:�vmo�i�?3��(��ϹAf]��B�|��-=�dc,�� G��+�*���TJ�53M��Z�9�&B�V'�r$<��ڐo��JRe���M�F���E?O��/fћ!5��fW�������9nP*e�U��"����6;��Ђ�2U`V�Z{�i ��4��g��У�/^� �� �{J��M�y8���^��͗;�B�L��}P�5ڊ�� Ņ.�e�T�2�5ຜ��YJ� 9l��L�de=h�]�����rt��g(4�@���.���4|��ϻb
�ax !�Y]����T؞)K������K_�g6�^�G����4W�6����wA�(��#�)[���g������z�a�M���U�*ӵ�?���Q�AP��|��|�P,�m�s�Ű���'�Vj�l4� �x懟T,#��+F��L��O����^�!1,������ɲ9"Iw�O�����9����Ui��t��@���m���S��k:sOTc7*8��}��v���u�����zi����Q"o9�=4>T蕬b{V���?�ԠP�����q�O��\n2��?w��f���+�-�=����p׭ �~���
/�k��A��ݱ���2�r�ǟp^ԨK{�Sô��8�
D��fX>x�>;{��0b�r2ܡ��`\���5I+莾��������֟4=���L�E[�E'w?�V/�"}�$H�V�؊�O���l~.�a��2VӍ�s����ኗ
E KG�v݆Fge!�n̿,d�,�y��o���ꑋY��k�]S��8����&�xg�W��WCG�v�42�Z��SC�����	
ڱ�d��u�uiN^�]��L�)������ኙ1̠��u�- ��9����,̸M��bb���ݭ��[�ڹ�p�^���������rٿ"JO?�^u�!����|��G�;���.~.7�r��OR�X.*���c[��*�	���?�,�M���wB�g5���Tf���z���sv�����Vπ���H����_����.�gF\f2�.�0pz˨.�|� �z�^:f��Z (��i�E�j����!G-3x��c��9Q[���kz�<�9�Ӿ�З����,'�Gtq=J�S��c|]�����Y ���;��?|�����$��p�cL�ԅ}8Y����I�B�^@S�:(ߥ��E �k��$�۽�{�E>����B��\P��ڑ�D���g�	踄X��%�!�h�2+� ��%��s�� �X�4��ZaUl {ST�,��C����br%[��z�nG�O �[Ԧj�.<B%:�����%�t�ѭ�5K��Ǘ<3�К���,����fE�ui�����"..<9e��[c�4��u^;�ȅ�+{�[7�KH>�QLt�l��lV�+�@/@����+�F�JA����9P��Ũ�֢9�k��d�(����)��i�G�� ��G�9`�Wt~�͓Z�E���H�\��!����~�Y��*�`$���ʡLY��2��[3�u�X�,П+B&<�VG�����O�s�?�����z��1��۳g�f����wb}G�eM���kқy^X�>��Ӣf��(�\{�sy,��6vT+���v?��*)�,?W�h�^�8ُ���$ ��o��-6�2�g��%*�jo��63;Vcv�����w#h),���ؗN��Ɖ���������`�{�9��2�
������OW6H�;N�\ u�tZ�Y������)��j�%��D��u��7,�_S[@ݪ9�`�.g=��=�H��U��k��B�/̊�K���"!���@�M�� �ޛE��-�ܭvl��Z_\HcP Q��R���~�S�-�r�_��Ujm=�.n�/��'����#т��/���������nra�=��z����b�h�@7��ܕG�.Ztb.lV�\��J����܎��~$�l�b�yV�ʎ�Zb:<��~��z!���K���B��y��	��7m:Xس>Oڒw+�ж��J��w��C��E	[SS:�<T-�U�����a��>�X�G�v
�h1�����쇊�"�!k�N�g��N�>RYX�'�W���|;��`>fӯ�p�W!��R��r3���$_��Ix*�X�ey���㉢xV�ݝ��%RO�~��"�&�w��<��gV��=�D��W�/R�:��������vB�|��3���~Pn휋/�a�g�O�a�LN���m�F�)��`Y*�R�ߝ�0�:���{��#��d:*,I���_�uP�n�'�}��f��Cy���+��no+~�'r�z���1ܫ�|$q5�$D}�U���)]��;���:!H��?�^7:e�tV�9�ś&>�$�\��&�2u�4	�R���K����v�7~�ڐ�����6~o�����$�Fp�aU�q���V�i{��;S������*���!u{��[��s;��j�c�d	��f��V�&[5���:� -���ocF��,��
�����}4�K�(X�f���-(�����W��V����57+|��~�U�|3�(��q3F�Ĵ���m[�G�0A�æ�x�����p��rč��;��_:3��t��p_�tj��?�x�+1i�7G��ޔ(��եy՘��?T��#��,i���l�!A#������8��B�o���?Җ_y���X�U�����p}�?��:,��{DAE�E@�AJRQ��.II��4�G�����Jb���$�`�y��<����xyy1g���}��^k�9@�}y7;Q4%��3�\d��{��_N�^���H�B���}YeX���A[�]峐'�|�`�Q�t� ~Om��.wP~���?��אv�T� ��;dږ,rDe���>�CN�A+?�y���si�,��%��n{<�9����%� �z��|�]s4�����ǝE>��a'4�w����@�b����H/�X����w�		��w��G��-�O�CK��9������8�8f��P��G͞���y��8�o����N\���C8!p)�XZ�f�r};��w�$������z�w�R�|�~����)Hv�����"��~[GGg8�pe�G�bz6h��_��q+�mY� �HA���?{�,
nE����;.�U�yrs��9D��U��>���T�Ĥ �,,��֨炵ۺU�}c��	��[<����FW;F��Eo��k�V�����՝��J���B �q��y�|�|S�D$ dθ��^���ɣFw�ݧ#�n�ē`�.����_ 	DO���K`�ɾQ�n�U��.$�|�:>B�d'bE�y��6���� ���m�W��v8���8/��D��]�`�Z�v�ی�:�f�?�6C��Z�YN�����
Џ�s0��s�Ah��}�� ʅ�ȩڋx2�4���홓x���ס"((�����Y����KST���(�� ���)������$��'�}�-�j爇�W�8pؗ�q��FvM�ģ, +�?�"�Lz{����%�漨�]���!Ga���^�D	�WeO��Ou{a��"���*��98t��!HV�exwP�k1�޿�y�~�N��YKE�D�����{b����E0C��r.wb�;�_�z=��o+�����J D�����R��r�
ѯ�Kɔ���,Ѐ�M�,��Fx5d�O��ѯ�zH��������l����R|<�V��+x�����Q�ӧ�������..[K���	��G�Y�@cQ7��2nm�+��ϧ���c��&v�:�����{��9.-�,SM����ҫW��h-�:�N�$;�3(k�������e��*�?�j��WZ7��(uHT�^��P����)�i������э�*=���K��/�rfڢ*���`uwO��)�7q�svW�'w�"'�9�DbwP��5Qk*���%*�$V��l��)f;��9{Jٳb��N�c&���,���I7�+��4s��p�b�cwm��E������)R�YςkJ��w���R�0��Ώֈ�xy]�C�@Z{ըw4n�7�����{����>���xS P8�}/"��wB6=ȇ�2�� )9��e:<����n�?C��\a�)w��� b�x��X���+���C��}��.����h����dw�;̡�F�����v��c��>��Κ�+��T��2�_5Y�:jE������Zj;�Alnr)�^x������[2{}r^e�[���1y��^�%�D#1��p���'�4��o��NI),�I����iHx�̸����6H���2�"���>���c��=S�����j��eW����e��0K.���"�:Wٓ�M���J,���1V�8�l��:�<4�@S`���s7���ZNlPKK��5�3;��!����g��ޗ_l-W�	��e�-�Dॖ�N6,��o|{���d�<�"���k��@r�����ƁCbخ��|�T1&��UN�7T%�Zak��VX�BBO�1��3�x��'����Y b\�@3�()鮑e�����N�Q��Z
��(��jCYWp�R�Oi�����;u�[�	[��$�K����$px:SH^��
U�Jt��{ �@2�Z�Y��3k�~JH��H�_h*#��xm��)���&�7���f����V$�U�
xl��y���WM��+=C��+�����ѸO��cw%��0GNw݀`�w|���|quS��`�'5�E���]vW��ĩ�	�K��̉IT���e��w,O`��,cG�����xKH;�x�W~]����P�}8����p����C�~o^�vnع���5
��2�Z�=ѵ��v����>��}v�1�L����q����sj�!.mΫM���/�S�J�����{U��0Z��g2ҙ�$jf%P/�%VP���O��8+��w��L�MX���8��w�A����aQ������5�C}�wJ����CTbי( �m�����Y�%��e��r���;��F3�$��EA�-�/�E7N@���&�]M(�C�E�"j�X�#��_Q�׆�x�"73Q>�%	���Z9�����sG���Y�1�9�wx�-���w<���-XOXVơa?�w�
1�e��+VA�49O{�#~�J�b�	��>�1��ןg*�������@��g]_�����L`��֔N���(�(�*�'�i<�3?�<�bp�EII��.>I��3���l5S��	œތQ���[fD}U�f��x/|Z�<ۢH�쇈�v�����\WU�2���qy'_Ֆ�Q�O#ݼTf�h;��a&A�x��Z�е�_�W<��h��]�7��&,�o�-�.��g]AA���ݼ��),�m��9c2�9������lP�f�I�y�w+�d�zr����0㗞������=�����Ft$��R�/�DC����Ą���7��jj;�����~g����xcj�7,��r>Np���9ahdc9 k���^xچb{n�c�O䔂N��	�p�ݨ�:bG�MA�bR&�B︗�[�5:�/�)�\�d*Y�'�{`�:F?8��S�P�e��V��V��\/�]#Ǣ�>����/���_��-�bf�����7�"R�I;]����Q
~c2��;���)�t��J�B��]bV��.�(|��<e��2fw�T8b/39� g�Aby��E�a�u\�2v9}8�8�����~��FY5�h�0�w Ȩ��+�A���51���J��ϓt�Z�;p�P_��b"��j���?�1���/��2����:9u����U�?]5��YTFu�mq���x�[��~^Z���X�����J�M�Z��]A��ԲL��5F4���Y��W5�!cq�,rq^�>�������3K�A�χ�jČO�u�\f����t�ݘ�Z�����>���QSY��W���N��գ�Cp!���dC��� *M
�X�P���XeKdP?Z��1P��CQ\�zG�lN���
~�ʯ˧�&�-��=)�m��%� �An=��������˲�w8Me	�����Hs+�o�V��*´�486ۀ70v}��g;fџq�Ӱ����f�)Gwj�`�խz��8R�gh>}S�KC�g�</d�
;S�����䯏��e+��'"��R�����,�e�bK�v�-PU���:�I���V�i���i��n� ���J��K�}�����\O��9�Y�^8l=`|&���_%�]��j��v�\�o�s�F#&�����0�g��@�����}=��w`�R�S�p��� ����?b��Io�])���Z�N�׊���`���sr��}
'yg�;�ٸ�\ʅ�.�
{W�Ϫx�H��07�v��%G�w����]��@"�R���+6�S4���\�<X��<PռB��N�TV�Jp�$�$=�P_?�q�9mɷ�N��}�����q$`.����un�}UG$�sGSՠ7O��A$y+^�K���\�~�|K��_��9��>M�:{���͂Ad��M��2O����Y\�������5�$��АW�/K���w�J��3��{�l��*4A{�|����^fS\��ɳuȬD��&���0��^����Y���M�	�Zf�������,g
Ҹid�;u,��'M~�p\a���D��v�!��k�X�9j'����D||Ӎ��x���Sq\�1G4�尠�Gʘq�mX�q�Cx�+�s֨�^lR�<3��Ь�<Eqݝ���҆�~U
g��]k$+�#p�o��=ӼW�&�R5va�!/򉰌C&�↯������B�~�ă��;�`0����GyEu�
��6�`Wt�2���Ts�6�v'��=����ә@�"c�w��쌺Ys*%�)A�L���!�7�0b�z��-�-2x���W���Xe�0ԉ�Ɉc�}��z?���G}w%%
{��/R�A��9� %:��j�����M��g��Q\)R�Mb�ų�]�aY�qT!��Ƅ�2<"W
q����%�WM����8��j�8��UvÛ�DA���*/���	�XA�홣h�z��Ԟ5n����ƔI��ry��<�i .μ�|���}֫0 ��I(���!b�<s����J��`���(�ӿ>U}a<j+1�s$$��#��Ӻ,4��߅}�[аע}��f�`��s}�6��;��M�3��$<�Б >�OQ_�y�Zԏl{��{�z�����
��9}9v��%+M$���p���E/����N��N��kL�C��H�Гn<cX�\���/�L�����O�Y8�pA�X�wp��~H-���\����pض,q�/'A�:�����V��5��:O�u�vG��8b�綦6{����R���w5I��<����l�j�ɧg�R��P~8����V����/e��t���w3p5u�@�g�ӡ�9�@,{��>.�I�����;{����"�Z�?��/s��@('���K�h �8w�K��)�-�`�uw8���"^	e[%~�W���q�(��\i�	�J�L}O�34�oPk{�;oࢴ��zN���We-����Т��S���%�¡�{)΅�ӧ�45�֩�҇�@��'�����]0�{-f}���>�:��}y��5i3�<O����a���rx:0���w׏��D���I��<�o��-��ځ*�lo��0����� ijz}��(�R�ng��d����$f�(���浑gf���;ļ��	+1�_=X��8Jb~���/Sf+Z��-z%�(�~,��ܓ�n��V��y��N�:�"���K����vW�C86#ޜ�a����`d��f�o̵��X34�g�JM��<�=1:��<��'"��jC��.����6�;[kyu���A5T�&�f��3K�$�:�<���~ؓ�a����F0�v�����)��~K�SV]k��@��s�: �'��qB�L��R�)�eII���נ�vKbȏ3!Rqhqw��sU��^����ZyI�\�k��,w���s}�v��5^ޛ+�Z}��q$
l�FL�U������
�sP�5w� �@ �fd��Uc��0O�/���Yh`�1����b'�n���=Ą�_2ߎ.�ogbFy���k��k����F�p+U��qy��m��m5v�=[S.U�%w���g�4��㋪v�P���}V����A��l��y��q|�}� �~����)fq�&)��?bbV��H�)*�v�	$Qp�yRC�k>,��q�ȴ�CnH�t�D�袡-�ӫ�Wi=�3U��$<}�'�J7dO��s:����T��j��� ����>81+����i��S\O6�;�BBE���3��g�C��ߒ����։<�{M%���*�@���O�6�E��|�Xp�z�i��4��x^��T���43ZZs1�}lD�>�K��~#��)�%v)�W�j�㇘`�
�TX���1�c����G���}wR��wܷ���ǄF�ϷX����r	l�8Ծ���78`�A�柚�i\�,wAW�vKH��M���͐��B}�.v�c�ԙ��7�+_����s��@�=	n=�d ����.y�V$�ׯ:�S�L���=6�N+Z�A�󘔔%���%[ِ��ND�,�(��f^���bgC�}|��W�<<$@>>�sU�Z�A�z���F��c-9�9d��m~g�^������Ξ���e6�s��}��0��EF�Y%�a*�� Y̛�{�rE-sn�{J+EI���k�AH��&�F(8�Dr�I�YX��ry��h_��k|5�ס����ָv�_��9̲̔?ix��]w��Ꮾ��K�^�A�ё�l���b�ui�'}�c�ʲ�������,y��A��������w`\�<`ld�G���NJA���7B�5^����Cc��([�޷�458}����:)-k��`��qGb]8�ɻ�2�6�5��
u��]�|�-T9M�w�m����^mT�ij�L.w��W}=��(3�@�X&k�hZ�Ϳk�og��4))(�(>`�&�z��Vj>C�x��~؛�5�a��\�d=/
2=�ʳ��ۆu9gS��\��R�z<�3ē0:{K����R��X�e�$
��>��Ii��b��X�_�0���Jӛ��{25##ug��4=�?:�XgG|�Av�kp�Khjn)�/�/������D��*Z��F��H3+��6�^��]�ޢ��%{u�%�l�%myM��c��K�h����w�C�����^�m��r�I|q��f�7�
�r�~F���;wB)|6z��-`KfS��õ��ʒy�n+s�����.^QZd��춓E�Y��WT��G�h��r\z��h�_1
@A-��އSW�\/ }������	2_�e�Tfi����n2���v�b)�Îu;u��.����r��v���Aibۻ�=�t�}�P���ۯU�K'�|m�)�:n�q�ʬi��Q�P3��R�I�7o����E��a��-���2VG�������q�)3��$��F�b���J��5̐��UTvTV8�Ȟ�:8���П��7��=�|�C�տK�,���X�k%��5�X\Y�y��;uqN۞��Sx&�+p��o��Lo�0lMLJ�` �ԘvǑ����`H�_�ў�f(ΰ���#��x�ksV>$d�ͽ㞰��JQV��#Z6�C_T_�|�  �T:H'mpl�m�]��u���Qѕ���C=�g�6����}�3i߻Uֽ� ��^�w�d��B����$��x\^���v4��26��_;qfk1��ˇ�7��W��t���,�gZ���ΕTf$�r�V8�ĔHoo@�/�-]�FS$1���#��.�a�/N-t���ר�_gnn����`1�{XB�{�H��cԡɤ6��
z�e`Э�bt���4|�#>��&��M��ZR���#�$5��Z���YB���A���b�7d!��^P����pe�`��m`o���ߊ��;Il��N���Գ�����ڗ���öRQ
�^x*���fb=���Ԝd@JT��	��#A��c�as�X��QzWG��v%���z��d��U�ڟh�H�|��h�M:�L[V������_珗{�o}+���BL�YS�_�̙��.�F�!S����N\���@,FD��K��{e%�&+�be�q�[��2mS��Qx:�)��Y"�@�D��k���-[�|�"�C����4��C�AC�)�[��<Ej���������	�,22[n|�
���)��[*/ {��O��MA�pm�e-��q[b1w�z��P��k����!�y�^[JZ�&e�l84`$�@����|z�~N�IH���.�w:�Ƃ
�;��JA'��ꩃ\���)���"g��<�ge�x�&�ֽ��&�D&�./��o�6��E^������gM�8���hA*��Q���͑r.�G�6b*	�
�X�$b�RC�<��#��B�W�]��N .T����xM��fߦ�c��J�:V���:띞���M��(�$�m�C�^�{Bi�I���>��q���7oj��*�;�vwo��^�h���6���v�Pt:��x��1��W���AQ�b�@�[n�C�^M���Ҿjj�4��d����^u�6:�8�E4+�����N��Ó/G�1�gUC�bbp?�e8��R��~�J����#�T�sv���Af�Hsy�{�>��Z���������}���o�[O�{�Bng�@��ᔡ߅q����?ȉY�+��B{3�����7J2?ɚz�����M�>r���׫̭���U���RD��kl�˭��'�XU�UWΫv+x|~$)�VOl9��R��Sw[��]�S �Z��XϥãI��n���"�;�U�P{�
'' ��M$��7_`�(�Փ��M/�;3%�eq�c����}x��j�A��p��ҏ��X���م�R0����P��.y��w!ZL�\�9IM�#M٫�7y���\�����N��YZpK\�����4%Z��>"�DrI�|yW�� �i�a�ŶNV��;:���է�
�a8Vi'b�QY�^Y���(I���lLW�9z�X�Ծ��r�ۣ��3xѴBP���JK��+f���5]�c�v�ݑ�]���W�F����R�X�%�0"�M:)vv�����#"�6��*vm���N�����ط�x|x�>�W��싦����/���9�+�����g<e�8ȂG��,��	����X!l������� �e�ݜ.a��NQe��s�����6&e�u� ;����A�{>�� H�=�֧������K�A��-#b0\';}��g�8<������p�*�;��O_��kW�K� ���7=r}N�EM��51��L��NYD�<+�|�.� ��V�J���>��0�:���R��1��ۓle��X���hkda�b|T��[�Pw�M�?�������xqj� B�cH�/ՠR��ZsߌYR�g,�斖�������ɑ�#����J.��҅w��
�����֞nJW�u��\׽�(A���½pF=G$#��D�����.Wt)[�aW
w�~��(ߜx����{T_iڮT؎�_�y���J�F�����|C����Q+}��
�ز}v��<��[�KK1�4}rvI���cC{��O�dq�C�>�h������V�xEݘ�|������#���('�P%�`WEUo2�p��Q�䴍U�/N:Npb�@�
sԻʭ���4��	��&/ ������ߋ��������t7��$��(G���W7��yH��x#�q"pKe"�%��'j5_��ks�'���D<6	}L�:.`�GP��5��.JJy@C��ᖤ�O����� �<5#�ظ�k�Z��5��Z���2[���d�DWyW�U���;�;QR���x��^�`�(�l��^��d�ڟ%���Y�@��რ˴��@Ա�Y�ch�tJ�x�R�R7zrjs������u���K��q�N�\i۱nq�S�(a�d�i]���4��Cv�?ޮY��bd8�L
Q����Ȃ�Ȯ������_%�ϝ�/�Q�\f��{�
�U��՞*y��f��a�6�@F%������U�D1os�+���R��E=��{�G9���+�lA5�z�ѱ�D���)Xtl�+xCQ�h|؝̹>f�Ha�O`��(/��Zg�66GZ%�&���~��
M`
Bed�b����MΔ�a����`qA �g+*�-�ndx�_~�����.3e���;o�������k2����p�	��>�2P�9V)�����-	��O,������Sz��i}�P|���ze��[wY4��mg7�C(�J���{�3�- C(a@qʫg�����;���3�V�N�*����Z���_tn�^e��'��~�����@ӥ"����ROv���Mi�g��#�����
jNO�����l�����b���7" AB����m����P0�(1|ېK��Rc{���a?�kܙ��t�_7�_5.�'���"�1!>>Z�N��"����G���+�<�[v���
��.����ևd]����+���	�Y~Xz�F|��S�Y���;�k�]45�qC�O��a3Ϗxy����dd��t��Ź�����L������ԅ|Gu����B'6W��.��j���t��h�i��a�U�����r��McuMs
u- jt����Ԍ�x@�y_'��;��YM0OO.������Q1c���E�V�>�? Қ3{8�"�8����L�ݿ0�J� ����HF�D�}�A�"�L��,������bQx�NO5m��?��q��x��ho]�;������ ���`����i�f�GwK��O�uV����ڲ}^ъZ�>2��W��Hu�`j����?�������uU&u���u�cBB	v�	��s�^ɜ*��!�y��b����#�ü5��ޠ����W}49j�It>��$ޟ�4����	Go�\��t����~���P���0n�|�n�*����Qp�٭�Ƒ˺��=�1�&Y��{�	k-�X�����H�o�-�e���diHAD�9^�8;O��һ�W�3y��*Pc9��iN�&NN^��.�'쾉�Xp�r�yK�'�S�_�n�:L��P!��#�(%w4�)jf����҉����Lz�d%Έ�6KT����y��I��A�௓]��NF��?T�)���o��bwM�	eXc3D�v?kc��������	�xpQ�||�� k�4H��h���{���I��Pcr��C��tֶV��n�=�W.��8,H@O�;�z�#�F��'}��@�dM{֧O 8�ө}��GB��|��*5�iI�u�B+K�ЦW��T�֐��d��)�i@��u����ǽ{�%���XL��;V}���OuI4#|f�b���G�T�7<���`������+��#�N�x)�������1�B����".����Zy�6�/Ga8�؟�f���f
�-�E�0�o�<R�w��ɝ��u����C������S%BUmJ`ؼs�X/Ǹ�<�verw�9��-H�P�|Ҋ��M�/@�S�{|�(@~�I�m�QI�M���Hy2�¨n���ʠ���(����E����'�*$����c�"�G�tw����e6C�%v)�oޔqj=���>p3����hJ�B�T�qH�� �����w2QX0~B�ˋ���j(�LJ�&��xE�i1OE)�;XG�i��C�_�H���5���%7߅�|D&� �jʜ�s�V�s1.2��#�O��l��:Y��#)X�ۏ����^�l�7 ܵ�����	�ZKsL��("��+|�t���e7�=^������L��z>��<���&����+��Nzk.;�e�:�^=�^I�˩5� >��4(O��{5���7��{%r�<EP��U��3o3��~��+��h.+�r
"��e	5�|
��5*҉��O;�Y�,ߓ��z�o���|Vjd�����o_�пc�^��,O��75��"`n��gz[�N��Q.{�@Z�Ίԍ=,b2��2��9CD�m�s���ط�˙���Ͻ��{��뵡���O��"�j�?����|F���Z�]�Vj|G8}�C�?�y�~0�����urpȣ�<��=Gz�Ma�r��ɚ� �4.a��&�C�_e���e/󱐌�_��,*�ɷ��Fx�F�J6bP,`��c���Uu T�(�[)V ��e�^����&�9�Up���7
��&JJr�9���Mp;�=G����Uq�v��eR�e771��b����i��
[��W�߫�?��i�6<lh��"��߻���w��a����h�	M[a�� q`��L6�ɯ�T)�����$c��$�X��#�`rR	���n
���G��ϓ�{�j����������񝇊�o�k��~�tY�*�	t�h&/;;4;Oz	R�,J�Jk����*3]LM��[iC#��}�F���`�aќ�����l�-�;�r\�bY�mn���b�w�H�*�b��f���VE~�6�s��R3T����PA{q��䪤�.�6���ꋶ+��M*�A$�=� %��#T�r[1�>ة��A��������ڍW�%��b�Q5�ggζ��[GT��%���M���h��q	�]��;PZfX�b�J[G	aW�Ԗ�A���6K��u	T���^��K����HI��!9�Ւ	�2Ȱ8U�}��jzdԢ���*.��nu���:���b�Ǯ��s�H�sn���#A����1"��wG~�7[i�2��p�]\��q�����e��wQ�R"��<�.�Y7��i� &�Z=��cz�a�$�J�n��f4�jCb#�ʽ���J{<'?��ԙ�D��#��Cu@��
c���5�� 6L]}�
��ǹqQ���|Pp���O Z�d�z0�����Vv�dem�q�+�Z�v-)V'Q��\g!?}��L�Z�t���~ ֽ���y�H''÷�k>�,T
��B�Y�MIR�����x����gAzca �����h{ �k�mR�H�IL�>�>�03�NɃ@B$�Zr!u�|�oJ��ϲ�z���Z�O֪�ZQ���=������SW��EObi�0bin�DD���'�x�+~Xӻ���{�'	�M>��b��"�����r���o�.����� ����7�V-F��,l�1����}g�6i;/�!ˍ�B�7�#Q_Qђ9�Ŀ��bN�Q����P׽�^�vo5p^�� ����M�������@p�"�)�߮7�=UO��*/a,z#muRu�5ϝ>��?Sb���ls�<�W��g
�(!W>N�R������3�u$-l_�:�D�F�p|dļ�e�7 <��B`��C�7�և7�'�駝���c������N~�<n���T��)nv"*��q��`�p����1�� 
A�E�X�Fj�E/�;�X���>c�)�e�h�nfθ,�gH�-��@�UyVY��� �����z�njKݡ��� [����q�~M^^]�7��/�<�㒖��&����
X�A��
% �a�#"6Y�����|[����7r�gβ��V?��F���ǥ�5MG��/��7��%����'%���|�EE�����v�� ��x��S2�ps�O�&�n�����;Q+�ݪ����r�؂�z�\����)9�d�|�kd��[���o���M5�y��hZ(mU�{���"���Vod%����`t�E��'eH�J��v����G�h�E3y�$Z��i�N
b��n�.;��̟>���PU�k&�ل�	�+���c�}??�˗��?�t�1鍾"�mm�������;�P ������
ğ��j���(C�:����J	�0��$P�\��t����ԙXV�q��뫂l���t�̿�v�tm�<���u�ģ�/)�����l�C��d�s�؀Q�mhi	�,h[+"�}��ң='�[��-���u��#���K���dL����j|X����� o�
'�7ߑq�o���<���A��\�aaDS+Z��=n)W��������J�b���U]��fH������~Csj�_�Z�nɯ�̓�}�HFG��h�'�n��w�DZSg�̈́�I��3�s�D���D��Y�v_r-���ȍ_��@�F�xn|h2���f�)Ĕ�k���S�m�ҬFIR��2�Kj�	$�CL�Y,��M(Ɇ���q�Op>��QH$'%大�����������KH{�l�i�����dm���M�t����b�*�u`�o���(��N�L+�O��u�A9X�9�B�11�d�1ƞ�ᰬ�
9�� �B�0��қ����X�X9�������Ⴙ؏�ۻ��b#�&VVb'�8gS�Ft[�x̾a�H������Jg辱o3ԁZ�_��%^n���N 2��j0�}�G����Q��]�u�Ժ��X�?�?�>&iFAäG��[�B`*d�i�����DKγy	ʎ��.�2����(*�ԧ_��aa���%>��/٩�8}RL�HK$dBY�!Q�j�1�:o[G�X\o௬��k�{������_5[����xB�	���]�T�#uQ��7��
9Z����QRǲϒ!T�7��Q�&6�o@w���(�z_�����=�Y/k��U����h{&(�^�;qI)c��܀��_T�p*R���`�����3yu�BuW��CBy� �'�eO�>$$�1�:�]�C[��_^�t�~�6�O�*�rT�F����ńA���
���5̈��6�w���A�>��RD�(W'x����IxS�x�-J�HҾ��)C����)��닉�k{�T=&>7��`��N�)��O��9(�VW�>�>�O���7s�h��I�l-^D��=뉨�(�~:\_�z	2�����6`��oQ�>�����rH���tKȿċ+��&���ƍ>��=���[��S�W�@�7�et������wΊ�p���>a!�0 5Z~�޷�Y'�$��`J��K/�����}n�R��6.��q�<|гU&�d���� �f�Ρ�F	p&��j��e�*��t'�d��_[��嗻C��H��"̃3T�u;���i�M8�B,��:��ji@�qn��b-�bq4F�Gl�kD����&'5tR�й�?T����9P1���܎���	ed��V4(5�[8��U�s�t�&��Y5�������@3]���;��U�V��zw��@��!Q\Y���q�?��޹/(�
4�<Mn��:1��0�oϳ���Q؆�������M{�F	ѣ �����ɣ`[d��.�ڂ0�l	)��ި�s���ūu&������a���r�I$�q����'�h5~��&��¨.8>�Jc���a�'�oE2#j�����"#S�ܜ�4JW���y�a�j����2eU����1<.J�8q�]�~����YS������q3F��A(L'���:��Wb����kFt����=b~�#��C�%(VĻ���q��g�4^O!A��\(�}+�X� �c�m�-)�uY���l������t��g��9���'.S�b*����M2!��d�G=��x����)�[��� wj��=	T(sֆ��6�ͻ�2S��MS�~Kym�������5{|�hv�n����c��~el�kt���[���U2!JX����}�k\��B/�B;:�%fr����E����+E|��~}"��V89���yN�W�㢹q��p��i���Zf�O��J<㹤Iy�c ����t'/�7J�GQ������~�k�1���;�·�0�ww�JkIΉژ/��X�3��ߛi��F-͙!�>�����I�O�t�,"��i�2�?J&����y��.��_7
����Z��#*tǯ�n���d�+(.�>��W�ϱ�#��x����/x(5��e��N�L�؃Z�*��yTQF�^���+��d��c���t!?�؆!�����.��R��q3#c(�A�P}T���8�YÙ㭝}���u7�vw��X�OF֗D˯zRU]�J2�����	.�k�����7��d,܄��]B �7��q�4{<ݬ�X$>�9Ua�:�N�`N�K�Nx�_���&Į�f7nP.M��p���B����pJ��@���!M�� 	��9������d�h��`}p�xr�P�ռw����y��^�-D%q}����QRH�ӈ��z��C(�b�B/� �����p�r�=���g}f�M�{�9jp�R%'FW9h�@�DF>>��˽Pu������H���li��L�b3���*/�,=�{c'�ؽD-ë,"�cS]��^F�ֱ�|�+Ц��Ih2m�����y�����h���,�� �w^��(��r��B�fz�\�X��3�N�B^��dH�����!F��k��z�l�Ǆ��R�ﴌ��"��ja���U�_��}�Z0��͖0���Mc��˙^{o�j(��۵��А�GJ�6b��������*Q���E� &.��'u%���7���c؏�vv/�ɔ/�/�|�O��ws ��6갇x���՛�����d*�[��%�D�]u�]nnb�U���I���a���hz��D?���4�eܨ�YyɃ����OdˋriΪ ~��~�{��I�B4� �wE.�40�/����m���kܿ��S&Xw�F-��hKM�a<p��W"Ȧ^���"�}����1�ReT�B
�w��]h'>}������io�����"\�W���M��[�n�˅�l}��r�`�]��߹;�	,E��E�O<����\���Q�sC�ĺ"������_�l�fA�Un�qj��Uf��In�Q�� �U��WP0a��^�}<�p,s�V�	��QN�:��f1C�DV6̫W-����(+�,�������*��>s�W:ȉ���?\�I�� �j���NA�D��¼_���٨�-�TJ� 7w�L��jWey�Ue�D�g�d
~c�=M��8H�J`��o9����XF&Y�x�x'�he�㴾�;��"-��z����|R(}=JY�<O%�0�ׅ��m�V�� Z2Oy��^�ӸnZ����vQ�j���ǳ��=ߍ��p��?��r�t���ӝH��/::�7��6U�) �5�t0�fD4�p�{�N��h�P����Um���vV�0���}������])���5T��<.��XRL�wZ�l��^�ܻl�\<uu��hX�J@��aV&���9�ql���O�	\�:�vMM͚��@���䆸�t4xW��~5�{^��\Y�����X��l�LH�R�ꂡK�07_��$2��N�|��J��N�l0�t�Ib#��p�۵�o7��8Ml�y͟�b��z��VT�:�k!:q%��خr^��4q/�17�f����v�WB��#)&�ݡWj�/P|Ȫ�E�E�]��0���I������ʢ�0�_�h
<A����]�`�S��K!�V8uB?@^�����\Mڶy�m~^IHi��J
�����r�(�|fHt�5HR�,�	��Y'ʖ�$��ՓhS��9�ݹ�6��C�ψ��М�5���.��4#Z�L1��e�`�l5�r���C'��yB;�>׫�م*�s5~sH8N�b�W{�O(�ƿ��jD0����ݚ�c��׊e���t�k�������8��Q/�z��vRkk]�����7ߍ�/�&����Q�HY�x��J�g�Y
h���b��Y��s�5q_��7g� r��������(t5�|�@\/ �Y�o'�7e�s4h�'y�Fߛ��as]RXK����>o��B��k�"���2T�� ����/��t����P؎d��{IHx)�H��mYm�p��c���[ګ�sj���dnwP0�M���M
��<��¨�c���6�H���dm�Od�����kA.c�T�7o��x�p��E6N�Ş�)V�'x�E�p�����-����1l�a�t�.kS�ܦ���^�~�!��� d��L@�ߏm�c�R��^[�#����|�;֕�G˚Y�Ϗ��	�vP�GG��F�����O`���Ӕ�]�͓��NMO7����i-.�s��cǒ��^�@��{
!N����-)as��Ň� \ ���M�u����O0CF�)i�>_�Ul^ao�����Kl�*l�艤/�۶W����&�LT��O���n��Sx��YYw�{������7{�g�:\]��Qk�;L��=K!4�����5�[[����1�z�_��3K}S����Žá;��	�g��8Ǆ��_��/2�����ꨨ���CRJJ�")�-�(�݈t���3��"-!)� 9�    �� 9� C|g���~k}���z]�9{��y��y�~�9>�B�PE�/��~����B��z6=��[������YcAHZFPE+���m�3_���}/N��ɮ��G%FUY����͎Q̡��̈����GS
�7s�&Q�p�Є{�ڢ;p:�d�J����� ��U������>�V��ރ�eȢ����_fF`⧵����}�o�7&W�RF�s���8UJ"�e��yw�׳b�����i@�WL}�P�0���;��(2�8q"I�hR{��y��-t��P<m����BWUi���W$�����s_��-�}�<��jb�����Ź���\�h�OO
D�t���S�T���^S�W�eˁ��7jxnV�z�r������ؿ�m�k
%�=`�u@2���F~����aBʞ��7I�Nc���pP^�|F	����C�~���R[SWr|��3d�rN�.�J05�67w���R ��X����n���`����q���F���@�C��<�1Uk��?�|�ϓX1 ���M�7�=��k�\�o��>��r������M ��wk�0�����%��f=�pA_H#wO�p#����ވ�+k�(X�,O%%�p,��R_�c���׮vq�Q�Sc���*���x�x^��.�P%��41W�SE3���ƪ� �|V�|6�=��E&j$.����j�`a���z~�
��t��0l��))���x�Dk�T����k� M�ب�|{��<�	�%��J���&�~�H~u�{T�6�@F���u�c;Rgɮ�:i���Ղ���Ћ߼�pY��9o�o� ��Iɚn�UEg��Ǌ`�������f�����!I��T ��oë��bT0��b�Z�ݪ�}ӎ����s9�#klbB	w���d��y�'Qm�&)���/D훹�/���;*���k��w�0�����Վ\�.�k��.ڴ������ݥ*RB�<�@y�|`�����pa"�v��r��Y��������-X��I��z��m\�� �zgY9gJո#{�eE����*zi�G���:b����j�'!,i�p�K�8st)���.����H�-��E�� ?�9���r��x[ٺ���g>�l�k��t�u��O��l>�%|�W�j���lN�6�E�������i�i������K���c  ɞ��"�.�"{�Ȗ;�[���
����K8�/�����0ֶ��4j4<�M{;��)��# �Mb���~4�����`fe�nQZ�B�;�����:8�}^Q�[+b\.E��qN��k
��B����冣�\����-P��衽��r����B�:z.L�N����t���H�d���������#UN:>u����ą�=e]H����5�?7�p��Wa��`�r���R�Q�
;�x�L�SO��0BO��W�'�XXb��q~��#�~����`~Fێ�:m�.��T�*C�t
?��t6.�S��	���=��+#�q��F��`^�w��;�cj�s�;�`ȷj���֔��������oQ���o.椒��ZS���tL�9%u���_
�������<$�t&��)з ��yƯ�E��#7�j�0N#�sr�p��c�+����=*�Q��>��Rn�G���)�N��g�HY6S�Q��66lB��D�m�Kd&6)��'���YcaG\�~��A8�����9pu�5;��F.��j����w1�=L"��C���&cB��@��ZQ������-��$
"��y4��]�T`Y�����Zh��ځ�g�ô�LBɢ؄D��VY��r����y��w".�5x�1FUo�T|8�tLLrr|�zst`��1��SI��i���;��$^\^��� )R�C�%z��1U�&T&*�=�BW���6���k|T�l�Fn��
N�L�zg+��'�*ѝ���$<eB|�2�O����bK!�:Ĩ�WnOm=�����nɊ��5j�B~������v}ĈOt�vg�p�颫��iCa������0�3Ά���g	�џ��5~ĳ���7����t�"ID/M6��a$N�p�.��|��
Bl$���\1t$�L�!����	I�� b�{Z�>��ό�eX-�U��H���L����&8������	�<y����˅�S⻨����oڧ�t�� ����vt��#m}R���oB"�I�����{����JJc�ՁgV����|�O�%9m�q���8�k]f��Y"�
j>˰�ֲ�W$TV�*��^��)����I��b#��ސ�~�����Ol+���O���n~�L�74U���$�����ʫ���O�����|�*�[D��i�z��q�o�3���,c��#"O����/������vʖ+@�
bIket�������qZǙ���J��j8�j�-gF�Vl^(���ߗKJ)�t���]X؊�WJ, -��WѾwo�+��3s[lJL�z<>1n�1������gCw�tf�̆W�@����~I��t�_�nn��.辵� ���q�cĞ
�h�TQN��~�^4��x�}��S{�q��U����Q�U|ٱ��Wh��g}F�Zh�-����ܒv�Q��0�m|?�����g�Ʉ=9�͢��Nl���eˑ@�}����J;�~l�6qˋvdf� &4��J�+zä�S��ۻë��|���l��������u�$��%�����2����[����s��JDH�p�����Wǁ�ǧ�g2�)���% ����w�`*�5��j�*-����k����ӊ�?�lH��lU���ϐ����O�T�%����n}Ya�"a�#+�C�T�嫇�-`�،y��/�	g��X�1 "�,ʼPP����J����u�1�zd&u��]����95���Q�,�w��7/f��~'ݎ���b�a^���͒�.�>l^�n��Ȭ�fnO�E�z�A��2/<�	p���{EA蹌)Ɉ�c ɨ����O����k����/�*!�+XRĴ�'�NOFn�E=ÞbtC����ǘ���J�ts�5K�*�����CeR����XJEt(mgm��u}q�����Ug��
�;z�8N�9���{{Ka���>�ۺ��7|����d0D��HI�o�PM�N�M���]�L�o����Ѽ�nt�@{\I�'�Y�/�a��w�_E��Ȟ����_�B�5]�b���xf�h�;���Y��a���5ܴ�g��v5�'8���w�#��E-Y�	��WU�{��h�M���UQa��#5�F[����A�n�N���	F '����:����&�y��.\��0Hlr>�il^֮o�Wݒj��Lm�pf��n��A�U��d��שDad�2����Z�Jg��{ڣ���As0�;�zy�_���:�6���ɦ�5r|�B��#�<��$�m��&����K^�rYЌ�#�!y���f�Nɝ�tT�A\s�uּ�z	K����ȸ��ۉX�>�ӏLJ?�aS�P�j�&��^s�/��*�N��D6�w�v�]$��YŮ'G�����J�T^��)l�X�=2ʢ�u����*���VDm�	�{��gi���#+I�B���UE1���l�r�A���#w:['�ϼ�K�޾&��d������ϳ'������$��.{���/�}�9�C�S{�ZB�;g"�\�y��*����r1r�lC�@6��y�gX�����f�\)�q��ʹO�]%F�}|jW��1��ڒD�дZjY�`j���5����S�T}����ԀAU8�����?����΁3�=���w��W�j��sd)�7]��qT��b��HLJ�EE��}��I|�pÑ]'�b�_���.����PH�_�u{j׫"k}<��k8\})�'��U<p��������r�����(*��N�#�/�����th�*4n`���y	&,6��bVEa���$�u���w��N����ﯺT�2����w` a1"����������_ճ�,�=�t�1ޡr�=8��H�����t��Pj�N`�4�$��ǧү2�1�k���uS?cr�sw�ϫ�?�x��w��
"����~������z�Ycj��2/��)&2�'�
�'�L�Ʀ�����R�y��Z���3~��ձ��؈0�E[���8�֟���
����M��L�ݰ"s.�Ha�?̢�R/uNW�y�� ����Ͽd���t�n��6!�oRa�vR����\�Q�����9�n%�]w�Q�����M�Q�1m�
�1�-��5���ȿ�b�A���l_�F�ܵ���Q:u��n��o�Uc2�o�@Z�J�NB�����A�*��8���{8<�>��&�В�M��c��.?�B,g|߄�8,eN�}�X��X�?j������Ak~�o��a��"�X�{ ���`�������з���K_a�B��Rj�����f�yO$��; 
)VJy�C1�n��u���Rs� � ��ox���sb�u��E�b���ZC�O��N�{���22�)��,����(�~f��{Bʨ�M]6/Ɗ/�H쫐1��=�'K,��=���tv�q^���r�\, (�gIs�Ѩ�zF�eE���(B�ʖoV��P��HP��\w���-�r�6!�;8%���\Yg�g5:;���*��QD�$Dd ��@�,��l��[!����EIgf��ԝږMޝa,�0�/�в`V⊪ǽ��4�Yسb�z�+O�F��q���J�c�S.W�6���ΟL(�v��{ojwS�&m���F}{a���O�Ur$Ȟ�����E���1������%yr��1�����N�bN8�W^L$o�ǘT�����	�G�c�^Y��!!H3�Ca� �qz�|�W��o�+�;�U�:���w� l����͠{�����
 q�N{�q:����t�k��cf
"D依Ea��VU��z�	\ȑ�h1��1�ۻ�pnCja�_1�囱gO�G�L�<T���0q2�+�/9�V���$�$3�χ[]�7/y_�:F�FF�c�}d!/���z��r3}��vGg��z�ZA;r�Ǻ����[W�K5+^��zPT;鸬k��0������j��Y��l�c||�ar�:a�r����� VW���zaj��U2�̱
�=��|Ӭȼ�hb"�@�^�Fm�0��"��!��QR�bE�Mof�� ��l�5orB�W���6����I;�G�����zДx��
�{p�M���Xr��
�"u1C�]|Z��|9A�2�v���`�)1�-P.���	g�%K����g:X�ь�>,TU-˔������M�4[̭*�*,@2����ah�U�qؕc���ی�7&z�KiK��M<��8ڞE�t�=5H�E�|��d�0��y�-�W��s��{�6!�|��ˣ��� �p$����1 f�✦ �@J���J�����;*w�t�0T�=�wB�_�wڤ�I��7�R�z|>���� ǹ/���|�}�E�'t&5���l׏�������^^�x͇u�+l��U�y811��}�r
=��1���w�t-0TG<�7�9Ѓ���ic�`���>���S��`ⱖ$���u�Ԫ�0�xo��M��M*����^p�KH��;���{�L?�*���&q���h_)�V@�bǏ�2e�۸lc��K�Լk�[>[�>;m����9i0�r<j�K{U�6ѻ���bγ5�5�G�l5���ܤ��$� ��vh]��d��/��둪�� ��RXׇ읈��.��s�7�[��?��
M�ȍ���g��Aw�u�#�4�~g��Tk����>E�Ct�g�8G;�����c��x);�ɘ�������x��xV2Q�9�$u>(:��
��U� Y�NT�t~�r���F����@����H�@�^�_:���n9�;����L������ڈ�_��4�!o���KQ��|��しoUf!o�S����ӺeG�n����ӯH���t�����R;��QD�}��|��ba����/��#amȧ~�6�f���ӓq1ku��M��/�<MJ���:�.�Z��\s���͉��e�bַ���v�����H�g��n��ϲ��υk3J��#��`?������pw��.{XeTe1�zz�R��̢�@P�Jg��z�իN�\�b2Z��,�8�1_l�^�ϛ���wRBe�d�%��ѷRR�L���Ժ~�čǘ��x��kG��Q
�����+� ���8ʐ?/�M=)g���,<��@�Y��B��������r���ݶ�B&�Ю��WY��5ϳ�k�@-Կ�� r�N��bd�UN�Օ�c9e��>�U�S�M�G*�I�Ŏ����P/��k�䰟~8'$�:1��wRΫ���\\|���#�NkLo��������?;Sܬ�I)\ّ��Y����n��%����}�庡`
Z����S/��Qi��F_�z!�-�<�A˴wI�����s�S������l�6j�s����>��p&&
J3�W:M�$u�2�k-�cn�bO` �,���Sz�3�;�W-_�\�'6�i� ���x�s�F#�1�e3��:���y�s\1&M�`�Z�w|�n���m|{��ԗ�����P1O��N3��3�GR�Ľ���@�����1����ˏ���� <��AI�\m���b�}�K.�b�T�S��g���(;b�~~��>�;�����F��߶�����ep�MH����<j�l+5EI��{w�i�A�e���Qz���,�|(2_�0q��ycڌ'E[���+�U������{~��V_�u~L��(�]�+�����w�d����%���q'm��`�+^!q\���Գ�+��%*� ��Ə��/�N�Ο��i�=@gG9Gu� ��p]�5(�Z��Uߟ��©��é9�M��&i��g��3Ry/��w�f�v���[u�������A
����>	�]��+��g�|t#G�Tk�2�p��NQ5�_{��r8�H���=eװ��NՁ�23��q
�J���K�/�\=T[�!���T���tA��S6�bK$gr������J�y�b��F��k]�gj�
�o�d�#��HCcq�>��U��Ԑ�M��	
�������x��-m�|���^���kz�A�k�t��d���b
Bk��*������g���2~L%L��\����j����$�����H��!A�T�m�ϡ\[�z$L��J���\Tz�:Rc�����LƳ�+�lK�J ���3z�R(�>�,i�+\�SF��o�yD�\���=IZ�M)A�"V4�`~d�e=�Q�ŗ).�%������T_��Z�~�Z��d��"2�J��N�L�ю(��k����S� rașTy��R��z�l����Y*2AJd���tZ�(<[䓰G�i%�����N�N3�-p������]�@fD��l�ʣO|��v���� ܇����v�d��6����� �k��)���"��ba	�3�gr�Qҥ���1+���7�'�1z"YT$˾^
�ޗ�C��ֈ�77�%n;'���LHX�0�5����փ�#\��?2F��Ea�`�E<EE��8'���g�t���������|j�UCra�6�kNV���.S;/�#��'�������:���;�L����s�^h�b��ՕX���G����eϳ++�]Q�A��4@��	�:�ʟ)o���|H"�>m��A�I���,�^˖�[/���j8
�T"���/�|�$��͹��2ڏ�Y��Z?�;e��Qg��4�nT0�_%���w� Ỹ��u�Nc�%�^�r&Ϲ���i�|+�n^�G�)�&��b6�gԌ���Կ�7������9X~Ƌ�1�3ry�Mm��m��K��8O.�#�;n�4�tȇ]�:3.Nmߞ+x���� x�<��v&<�:����v�z�߁ؖk	��9�^]7�l�J\O;m��3�t7�;���vw�4�ţw�g[��7p�+���^�
<Co7ST�lix���$0Ya�(�F��X�D,<�S_��Uf�vA��i�B3�Po��H�/Z�����ŕ��-w��	,`��ԋ�J>.yfO3O�Y;y�zI��[0}گ�GU���^�80i*��[>*�/���+\� ����1P�l���ӥ������i��p���"ے6�П.����L�5]�t�� �6�<$n�)m�/c��)���G_���X�ߏ�w�:�=�m�d�'�.���������着D"��)h�<"�%���N��hh�Kq\.�ё��o�(�Z����䋞��mww�I�p��xֿw$`b'ӛ�6�o����4��t�Cb_5�j�F���N8A%=�h_p���5��-[V!��-Al3�ٍ+)��߆�gk�Qawvs�Bg~��'m��Mt������}�>�1�[0Zb@:00޸��p��d��ϲe� ������k?a9S��/��e&�����.>�)"�B�h{U�`e���k ��V��kk!��-�� M�Љ�cr �>%�z���o��j�����u��,��x��ͥ
�4J���n}v�v6/�ʎOw��,�u&� ��T�rd�;�	1�-������>��o$(��y�Vڨ@ޓϲ?����F��w\	r�{ LgMv0^��o5@ެ�\�����!*R��9�g�	��?LM	_3#�ƑKǧ#b�mz��y��ʀb�o�p�	=*�@����5/�c���ۓͥlS�	3�K.�7XS�ү�9���tTAhu,��lNԟR������n�;=Z���ÿ����R?��۫D�@�?bm� 966bB���aP���)E��_�!��f?[�X��{�S��e�u=7kB\��*�H�_%6�M����0���eS*�C@4�J�R����Q��B�1�9a��x ��i�
�ߡ�} MQ65E ���h��/��a��;����{�^"����΋�/㍅s��e9$	A�&�AM�UU����-|*<ch/��T~��K-����BoPT;D3'��O/vbq!��F�����M�BN/��Oo�O5��BG39v^Z<���������{<0��Lb �S���D�2��4NP�R��F�!$�j6%���R����<D�a����)5�Haӧ���?pvsT�M1�ФF=1U��B�5����ݣ����3(��HU��p
S�l�(�;o㎫�|�-�N��(��.����smT�NN����YK$[H�o>�m$��4A�C@+$��r��ﷀ80��44t$�wS&�����M7���Sl͔�k@��'�[�*O��0����6�G$D}�B���Ћ�^�����Ɲp�D�����4��$2z�W&��ZK����iX�G2<����%�!��m��@f�4����Ab�q?��6^��ז6 W��Hm�d�B�}�W{,�U�  W
�)�ץ��F���	�)H����C���DN�)���g~�
�n�r������K�zğ{V(�E�J+��[S$�;>�2ܤV�!��|�n�ǯu�20`��йR%�7O�J�<��vT������iEʷ[����gk�{
��<�{~�Ϯ�;�n���_]}��ߝ`L�W!ߧ����x� �L��yT��x�����w��n`�d]�U�r.���)k�tv��n��c�2ڏV� ��?�"5�6��:hŵ���q!��ԛQpp��
��[c�V9��G��cO���ߏ�ʎ0��[�ޫ�c}R�ȫ��Y_� F ���Ϫ���NA^�Թ��`�BtXA^�B�h����B��%����y�J�=��)쒱�r��"�[�9��1xt�r�wJ<�й��h�:���iW�p�9���YU�A����t��ªc�����?����p�Y�w���S�e��i��t���3�>�q��f�-8/q�����S�zl�.��"7�jEF��K��#��+��}�>ݜ9��t�6R�J�ݷ{�����Rqg�'w���@K�{.�@h��sr^�`aBf�&N~+(�[����P�����c�\��{12�H
��@�j7�������i_RO�)�̆y�=
��)��Y`��[{sO�(�O�X�%#F�6��آڟ.C@B��
��cMZ
��#3s|P���	8M���VXOʐ��^�;\�Ь�$�8�ͷ�"uʮh���z�>5�/��ه\~�e~_�q_����z���?��<PDۈ-��EvR'���\8}@���,n�_X���ߪ7`���m��v��/���n�ߴ�d)u�_�EU_D�����Y=��ˑ�X�c�u�}s��H�t<72�p��V�X�u���p9����9hu���� �M&�p|iȝ)o���`�Zտ�DR��`��Z8́v	�mkj+=r�q0�Y�<P��h��Ňp�m	��d,Q'�[SΈ�s�"��}I�����%�d����D��S�>�.F!ї�����'�\���@��p�̥�&A�GV�kkA�Ʒ�o����&$�I�H5^oo�ET��K4��q�7�nKmѓ-�n�p��8X9�k6��yi��h7w��?�i�ЙKy���Kr	��[Q�-��m�_�B��Fz}#������� ۫���A������ܕ��>�_RJhb�iȏ������VP{6J�+0/�__�O��f��Y������&���"��cw��I�>o��HШ�ۋ���Eɕ��H�j)��6*哤&ѵ�`/��1���):�y�yW�p9�����e6�z��GM��y��S�ͨ���,J�(7���[���ۿ�-�iͺ��V�BrU�G�VΝz ʴ�w+y�CZ}ՏQ�W��+��O�ߌ����CPQ1���D�3�aX�ۤΌ�Y���زd;ܠ$�(%
�92&n�e �OHv�tNT����r��h͐�ԓ��x�`_��P�Ḕ�1����*����` A�)>[z�#�g�#c	��^-+Z jd�,�� j5���L�H=A��]�'k@l[���a� roW�����н���i4"��Ƽ�g0.�w�&r��) �E#%��69o2��u�画0��-H4!}Ɯ[��L`��/���[p�ap�,�L�lX��b8#c����ZV�I��x��Q��Ol��Hl-�%$�_`�}���ܬ�X�y������硔ܾ��~W���c����'5��ӭXV��}���$�^��~��>�-$�=I�2.�Oy�^$ KE:OF��'ٵc �5��2�@܉ޏ�Ы�fm;�����T�mH$u�S�y�ү�S�|�Q!|-^�`Cb@.�O�~օQ�΅��\n�ն�!��� ~ H�����G_Z�/�,�^��M�3���#�g:S�WЋ�#�#gp���1)2��������`�Y�L!�����;��ͮv�ՙѮ��4���!�cD��Cy�h��/�E�a�L��b 9H�c!��=���n���e�юq��l)��5���������􏩃Ǻ���b3�@_���?i�������Z�xR�����R�w�>�c"���(�U.��푒&��.ZA�1qD��;
h-8�V�$�6!;�f��O[-�<-:�ͫ��\�g�ƒ�a�<]7	&X:����^<��{����{tBfq�eM0Ú땄f&*�TW�u�?� ��R��8�F���mL[�67t=�n��cN�����D����� �-yQ"8w+�y ��H7��^GN/�@&��emS�	r���J��mU��x�o������ ��o�s�W���	���qaP�c�� -Fn2��ꍚR;����ށޔ<j�W�4OL�HLZ
�������b�j�b�ni~ΰ�3���2�\l��l���[�J���۪C����H];�;��  ���AWװvWڗ����%�]|�3�����^�][T�v��7���_j�Q'�g.�3p����9��v ��;5��'����oIo���ؔ@�14��ǿ;B��i-O��ׯ����X���3��z�Й����]��p������$��3�^�{"|����j�[i�3?g��;���o*��"�م����U%%R������6�nc`x����IÌH�ו﷈wHpo%�O�@��Ҕ�� D�;V�.d�C�%��� ���dŗ���Q���f��7�<�6���ʣ��-�5��]P�jgD�K(�7�r*ͥ���z�}��zc�׌�����R����p�x�!AD�=���Y��r�Z�ٶ� ��г���"�32ğ���Y�j����)#� ����'��ک�#�G�x���~�!��]Q>�7L���̣J�`����:*�'��OM���-��çV�.8�#Y�Kϟ��[��_'m0�V&`���?j�,����ro�f3t�]��?dz�o�aO���Y�V±r��h�	�;�1p9�֜��%��&�()�e��?����.��j�+�"D����X���P�8|A�0%娆 ��#c5��%W�v�%���&gZ�+�H�q�� �e�[5��%I!������P>2gĜ-d6��1��C�;K�JsK4:��Oho_x�m����q��afv�#X�O�ٟ��m���U��)�I����Q�/��`o^e��y����5�\�������; �������P�E���Ku�ׂ�nхsa�t����0�ސJ>5f���.n�N�֐$ :��셈�*\��x���L8�Z`Ϛׇ��9��2ľ[{��<܇��2��07�:%��T��Y�G�fR��.��ES\���B�Qh툉��EI�痧���»���m!r0���R��iu�ϛ��q�@7�pd�q�ФQ@`&�j
!|��*j������Ǯ�����u�V����r̲<<��Hۚ8�O`��{t�#�85��/��ǉ�8��A����=_���1/׳pj�:O�� |s��o�d�.�^���77��&+Z���SJ�ƴ���J���N�W�R��z����''�O�X��P'A���n�۩�Z7��<^a��I���lU�����k:���*��Ȟ����P��=����Nj��GZ�A��cՀH8�=ݍ�QBb�Ao��L��cp�X��EY�.��=Ø�g>��O8���L��l�`�	���${BW�����Kw}D�kZ��<+]�Nυ���;]!["�Ϡ��B@��:�|聘xE���+)NA�r(�s�=58��1-[!�Ng���1 H�'��|)�M�����?�b����YSN�����1�vEx�sP.��sPZ��x������ssm�l����`������xr�o-8�<l�ɦ�}{W��LX�X�l,(9突:�o�6����#��kF�R�����q��"�r��2��	�h)!5�!�" Of�&y�� ���\���V����kd^z��h������A�OK&�B�x�k�A�%)���C�N:[���A�1}H)MG���z��X#K(<o�c�����ж������0qՉB�?�[^����@rYT��Gc)u�-3_η[%�F$=�����s7߹��զ�]��n���q�:�u��E&X��|ď�k��*��B��>8#[ջ�1&$$�;6�"�.a	���
2���kO��ft"��fe�~4MS�S{9j��;�����bn�J�M`9����r�}��#�+i.]�����>��KJ%4�ZJ�?C�1���QT��@��>�l3�~��!XO�o`
r���������Q������|d�2�x�����(�6��V��n?���
y9�F��"g����΁-x�q'�B�}��烳��C��HA�������F�z VAΥ[�4�#)�����at��@YT���������c����f�G��vD�b�����xI�`�[�4�i|��x�{�;����U������kC�Ho��FNj�������6@*�"y\��U�;��4��Z����i�g�N�oJ4	H5�"m�,MG/��^����^����v8��~4�s�tL\^ϔE@O=./p ��67����=���p!Gߞ�ҹ�z�N��Np�i�R�5��)�5���#�fC����uǅ4��ʈ;y��]��s�0\�n�܅Dbp�u
a����Op�9c�P�����@����p���⁹�K�Ƭ'NꍷF�����V��,i���X��`\��rj�;3�W]vU��*? ^=�����T�����F"�ޒv�z_����DrX?�>V�����5o���~�&p�����Aߺ�'R��p�"gL��gB�.o(��_i�<bM���F���B����]�]Ӯ���o�X1᫸�LD�V�+������R�__�wq�U]�I�2BB)+�{R�<�Μ��]�x]�H�nBm]�����{�ɮr�h����X��H��ľgƀ��<��,Ϛ���R!��+X��Y�d�9|eG���s�K>!ê��8
N�k��-�� Ζ�󭬞�����Q��1g	.�R�l�*��Z�U»��� ��a�&Xv_Y
���|��&Vĩ0O�Bg��Gf����GD�像�Boj8��8単4�J�͋��L��)����3�=��,Kd���=����_�m�Ʉ������H�_�"��:�p�y������c��{Gk:tՊ_ޞ�"�#��)����M�{V~HZ��׋X�Az,Hl��1c�߱���If�G�3C�t.Ժ�U$�7���͖(��ԈI���8��$��8f��ԗ��_�(��|~����e�OG�Eo$�e�A�̼�hs�&0f��pF\\k gq��t+	��J������0+wA��@�]��h�s/F��0a�8�2�R�-j�e�X����x�ѽ�	TnՐ��z��D���w.��rR��L-����@�ĳA�͆����o��]E�Y)��1��".�t%���c��4�b��0����4��8��"�rpvt$��'%��`������_�:��#�J��V.�nY�������N�q�?��L�7�P-I�`B`�N�:~l�,�F伡.����#�͠ �Ws�|``5幰�])��f��Ø���t�&u`�4S ���U�����}6�7��Ō����*�G���Ƿ�rᓭ)~V�'3 �"�F�0����Չ���@
70���~ȞJZ���j�${f/2V�xﲨX��j~d~��_�5ԭ��΃�@�;�^�#��|��bs����/�����B_r����;.h��v�����7�\��T�$Y��I�Ĳk�[����D;����2�N��ͳ� �u�՘gAg?R��t�̲?�/H����_}-�U郎�\���S���*��.�w�K�հ��쨣�ѷY� ���Nɱ��4}�b���~i-/�d�^�Qͣ�(uv��39E� �����5�6`�y�\���P���+�i����??	'�IP�M�����涚�eּ��,P��ޫ���?c����;�T������z�v� ����D�pך���x˙sy����mb��O�<��i��>j�	&�y�^�N�بgk���$�t��7r��J���\��\�յ��KK�
M�{33MPT�<>^���@�ۯp� ����%�vf[�)偝Ebb��o�ž�Vb��̏��W�\}�B&�'+�Bx�a���Ow�Ծ��o,�������M����G4���
ڝ�������_0G�����"��<�Q�w}g�Py��?�ž�h�sM�z� )\��<!l��B�װl>�z��PJ;\*r�ߋRk:?�����3��	Zm
{�7�1?����̱ٙ�ة�LtM��[?I�/h�W�jI���@�u�;�5Ew�z
�^�� ��S.}%M�6�)9�w��}��$����o΍F���LW�� �L�zń^z���P�q�⺵ԕ�+H�Ry���@�[>��Gv�L[�(�g��;q����?R�G
X�-zE!^>�K�������{�k�q����%e�1�4�Q��h�k�;��A�:�pb��l�8�8dH+UM�O{���8(��sb�G;b�N]�o�l���>�?]�[���]�I�(��Em ��i��G�\���uc#����U�F}�����b�i�Q�>	H҈ɅA����
*�O.<|�f����������8WZ����2s�^��ptzt��xؒ��/'cY��z�$���x��\�����嶐�G=u�A��)�����A���oȵ��5����]�7�
�.a!��X�N�I�{��t?�K�;;x�hg7}��2ᐺǸ��ׯ&�]�oG�Q7�v]�ŴG�%�U�i�{Vjp������xD��u�ErvR�Y�� `?AHid�,�� R�~�I]5� wEu)����^�u^I��V���RHFM��r�R_j_�-jyOW��U�k��W��+��5�=���X�l@����ۏ�1�J�C�o������a��l��d���l`�B�{-V+;�
��L��5��C�3愴����Q�W" L5EŽݘ��U��w�/�%�4_Y1��s%7ކ�R���0�I��^V�L�Cu{*�v� �g�+��w����3� !�� �c�n�r��
e�ـ]m��m�Kx�ir��Ŀ����%��`�#�@,�G�!��tEvYd�p'_2yh8�q�q�����HA�P�����tF]@zgΦ���g��&,��ס������2�i�t�L������mt���x��$n"CsO�e��!x��CWdU���C�Ψu+���u��%.��8�7m�i�4ҿ�g��<�)����l�o$�����K��a ]�����P��t�X��2��q���*S+��]���m7����S�&�'��8^��Q/��x�1<,S<�>T�5�^>�&J�k|̻�ru2����m<�2{�ǃ����mR�-���Gq�{ܼ�������z�޽�%4=[�[98�h��W4�����'����f���U�.O�%�6�4�56tL�}�n%� �̶����m�%2��筰3�uX=�$����k��iJ��H��ۏ����V�z������:�3)y���$^9��g�x���Q �3�;�3�#F��΍�f�4^�;5G��;k9%&�> y�#�h\����B��W�}N=tx��
ĩ�Dj���
qa��&���D�����aM�]�p\��Ea]�""J�^�G���ґ�Kh��(u�5�D@@@zOP�K�:��BK��L�}�x��}?���t23gN��}��Mfr��2�Tl��zΉ}^�S�j6�u2alr�2�X˕#��������L���'�t�@�n�ʀ���iq���@>Z9N@�3���6��h?'�Ӯ&a��H�O	����a|gO��\E����ʇ�q8X�9���*�R������ӐC�1ev�)����4�X�o�9�K	���!
+�WoO�l~"|:?p�s��Y�ȫJ�{�4��yz2+��^WA�
eQg���K�wE�V�Q7����sH�._-'��/ �^\�5�󹾯r��v�yN�>{��M����Ҍ1?Y��X��"2}[�~�ҭ=��t��f�D`a���՜��l.��-s\QY$�KJF�٢�ܲ7j�Y�����8���*��]��zz�.�yM����=����tqV�����v-���x�{6Z��ʗ�̝V}�A:�OfV��>yf�c��5Bz]jm:��ܹ��|k�Z㽫�n�� $>}"u����m�����pFf&�;6p�����Ȍ�{%�2�&8��!���a>������R�c�Jv6Jv�dg��Hֵ��d����3[U�`(�gȔ�����������fz�� Y�E���N<CS����=0���s��~���q��ʵ��Y?\i�u�w�*�8`溯8��`�K�M��ޭqT��᪡/�u&]l_A�X���e|Y_=i2Ns��i�������Hc<�n�t]��K�Z�3��9�;6��ǳ�'>��:χ�,+��ȶ0�~"2�8��:.��R-�2�Z�#��|��ҋ���+�o��6��l�>/�Ђ�w��,��}�A�@�!�xb���c0+$��:�8�Y���~����1�=-�V	���w����%u Yx{M<�2�j%W}�{:�1���d9��$ĕ�X#��²��:+��I���B�</8��Ռ����ȸ���y� r�O1��d��؜�L���fzg�~W��,݁>&�~z���#^�5G֐�[���#6{7]^N� ���w�Vp3�X��Tr�Oʫ����z�Z#95kē
0�镃�	?�78P�==��W��3us7�I�ە�Z��?qM�"_��H�O�e{�0f�t�bf�`f�����pn�����/E��?�e��z�I�f���wŗ�@:��N�r�H#�2�TJG�|X��R�O��!��@l�h8`�BL��e�vC��Yi�/޺y*n��)t-��₨G@�1�1r�������~�ͣ�1��n[��Vz��T&7 M�o�2fr2f��4O?��҃<��*k�j�D�Ʒ�_)�?�E����B�?m����z�x�TNn��i�N+p��%��m��X�>��B��`oq��T��l��F�nL�6��N�ʗ{�Én���_WۡBPg�����6i堾e�s��#e�Yj������E|�*m���4G��ϫ-��;�$�;p¯[����ٗT%���c�%��P"�"cNwbp��K�����(���E=��]8O\�������������嶟��K��b���.�7�����n�j޽k��Ok����������S��oz��jߛ6x��X@?���t��E9b�3��Ҏ�������S����� 4�}�]�7��B��A��6+�&�О�[��] 4��；��c�T���ESx�
��
{����Ș�Y�l�3�Uos���w:�^@";S�k�q�쾮@�X^dK�OAt�����]7�(Μ:����C
B��ʧM���)�a�����Y� ��
b�5�j�8�	�	�SW��C���� ��Z��^�b���•�L˽��S�N��'/ĝ8s{j�	�25z�O� ��3VR�������G���@J��:ޯ/g0Z�'�4��*܍)�`�EY�`��?3��-'�k7N�66�)�z�uQqϯ��"���2���ϳ.�}�d��e**EV��	� ��t* C�W�$a7R_<�#!Z��w��l\]I�g�	a����o�@J�X�vXLt��R~����n-k�_?w��K5X�_����c��>dx!�R/�qt���%��ޢ9crc��r��������ڧ�/Zj��|��"U�g����"�m�%Wֶ?�nw���x�v_��.@T��J�?�ܟC��:����3�ţ�|�Ej�F��#d[�孏�|N1���,�v���gw�l��!�<ǀA�[�=�9m3��Q;ϙ�G�f���u���A�|m���;=wý����3`�5��`#�qO6���_r7��}()��cOm'��NO|���?���U�滥fvZ��%�1���� �Al@�  J�����t�5o��V� �˕6p:���Ѽ���!��O!V]�jN9m�� 4m5S�FE���J�/�*���̖����n?���Q.��kk̛�~ԝ�H�Z�����b_N2�^엻�"#)Ȟ��p�˷��F��>�x��	�ష����u���R�(6O?��7��+�����L��Ypv��*/gcO�O�kU'�UY�����U���2ڂG�����K
�S�b��r ~��Y��u\l�~A(5]�퐡�[]n}Z�qʒ?��
i��`RN������_��i���,��yO��.�����=Y'��9ؕ53�n+sU�^�;��p2(���Ĺ��8�q�sF@����'W�d7;�#dw;U�r��i�Ͻ�erxa>$���9@���yOy>���ߡ�݆S��h^�hx@U����dV�R��H僘V}�t���ⱖ�8Ks���E^��Ԕ,r�7�0���|�W����2��F�������|8o��*��덻"�F���I�Ĺ�P�l�,/��:��S܈z	�̒t�×���\����9�d�5z����Լ;�q3��sť ۵�����8���ŝe��D6,�������|�Pw[��T��o56���khRGr�H4�m>`nJ��G)��`����:�M�;М/lʏ(�RQʻv�@{}�4Gs�9P菇�2:�I�ͨl	㙯G(��4����z��J�j��7X��{h(gF�[C?��8���������Y���![a�%sU�Y*���ʷZvf�oL�c���m����%6]��Ļ�d_ҟ1A����l�x��
'�p��V�KŴI҂#�-�u=���'��f��R�͜�]��6�2��.�;���w��
hFH���5�2����g<}���~x��#v��t[�K���~gR~�U�}/��/>+�}W�4�Y�u�y���5��*�@?�3��P�ZcՙW�`� v#@dn٦����ZԢ���.2�:yq4D�c���2Ax����Q��7P�ag=�Χyu~.�7�a�Q��Ө�]x{S��M�۩� 1�q�+ot?�Y��c��t'-�#������k�]S��
�ͶȬ�N��Mv��s��t�n��R��p<\@^\P��
��������a��������Vk�&��ai�]�H�5���[�f����L�$�� �xb��;���B6? C�r���L�~�hG
�"PZ�<���fo�Q��2�c8�2��D�)��X�����=I��vo^����S(K�[Ăm;09�M�Tr�<*�*�T{�� �|f���&��j^_w�|HY�c�j��Z�l"$t�D���j|@��~� ���'=��r4�b�.A�!��#x��1縦�\3.�#�R"]�����?(g`F�l�w�k��+e�c���olb2�B2	��"�שB��g���B�����$�Yce��|@������,)�\��G�w�zw�X�T��8����'¾8�H�}ac��o���cL^�)��F���|檝Y��r��G�V���ņ�[W-W]kO�.u��:y|<K-7���ty�Tw����`ݟV'ơ2<v=�w��PX��������(�^��q�ޚ�Y�����lRl>s:����Hb�g]3�bsn ��p#��f\zO�N�O�eo�0SH����;H.� �z �ƎeS�E1s"��2�~��e,qi���̞7z�����9/�����W���<,b��4g�	���R��Y7������3~�ц�h?Z�%��b|�m���$�� �����B�d���Dws��ak)�p[1�Mz|�J�Xi��=F\Z��^�.�!.͇��(��gԷ7������̾+8/^�k�q�(����]�U�TZ�S�l���PK����mȼ�$h�'�g����=�`��q*^����N��d����	}�;!���A�U�8ǘ6ǰ�:SY�W�=cf�{�]8i����@ePl*&ȇ��n`�J.vC
2�m0��(�hbcc;����2�?v�%J�i�'Ԏ����Vz��x�3VVl��f��Jn;�[��w�5BQQ���Ѹ�:�t,�~Oz��}
��͘����̀}�sY@�4�Q���$ �ݣ���-�!�1��i�J0bR�^�Ɩu�!u� ��=,s yI��49�"(Ή�ZtU�뫦��"�k�������� İ�A�W���D��_���mݜ0�z�{�9�G���� ������j��gj2�����l�j(�۵��� �P����̹[�܇F[W�.ܻ
��{-]�� .��MO&2D>�5��Z_-��>ӂ�vE���	/��|��"堬�Ƈ�v3��F)E��Q�L���F� dkvr��1A_�) �������'����X��@��p��'Ov���;/�1At=�-U,tk�� p��+��.l���`�"�2Z2֥�h��$�Ǿ%�����=���=�~y�?�̙��������%Ģ��@S���ӛ���>�J̚Ԛ�{f :Y������+�DiP���W���?���AAt���̲��4�C~��C�"�湛���ư����[͉�3�t�_-����ô��~��H�_�$��l�h���20K�A�&n nV%S�{��}6�t����SPTf��<���Z��I����@t�G�H�y��DC�GȬq�jď8���*t��D3�/gfg�i%�n�,��ک�w3G%�n���|([�f���^��9K6�[)����&�F!���\�N���V~x]cq%"3� �ڦ+�H�Ո�x�:#w���B��E,�,PW`��R�����^�᭍�l�X`��S[��'0>=�����f�I�����RĆ���u_Azgٞ��$����{i�[s�7{��17?�|��"����wF�!�������8���
M�W����:So�7Dǫ_�M�&<���eC�˳��lp���X��S~������Ia
�404��|7�1�KXR��TDD����0&�"��(/�X�qQ�Wm��u�!�0�;��
�2	�h8�\�� �lm��0�ww�S08�1XL=�a}U�;�S�뇭��9+���K��+��F^�����˗�{=�:�Lj�
����oЎ��N��z�����$ō�j�;�Vi\�qJdF��"�[����
�� {���EԚ|�[�ž[�	Ӿ.�G��n��KKp��,	~% t]�Ҹ}9i��L��b$��b���m�2|�@fв�v���5ZfJ�}����T�X���u���B.�fl��5�c�3�=\êӃ$!�Ǽ:
�;��T2z�W�~��RZ���{Q���C+��HhUV�jʲ�݄h�s��׋L��W���bh}FC�V2]�I��&�؋�nĨ�o�qpP�Ɋv��%��b��P�mu��Oܙp)�IrKr��SFG�q�[>���t��������0 ��9�����e�J��[�4^�\��0�c.�Q)�hoʥ�?661t����
"���4W���?��3�z�Cxnжp��܍��Q-��_u]����4s��w���10�v��՝<����@y�e�#LW�QgΪ�u����z�J5 )�g�޹���g�*S���I>�Q�N��C_z�3t�5��8}�|f��ጧTVM��=H� [�R�\w�g��_���Bޔ���G=_ג8�E�RZ�@0~�W���&�����~��d�I"<�su��_(sų�Ӿ��w��K��`�b�H$[�N�l*T��f9�͚=K{����
:ss�5�|��8K�r9#:�Z�����y_H�H���Տ��z��6�W��QJ��/`�Aν3F�B6/��� Wj��u�'��t��
���� r�S��MB�+�J������MJ�R��d� ؓȸ�\;{V-B$L�ӳW;?�EQ1s����	~�<Qq2�lrs�����3��3�[���q�,
(�����2Kog�����e�-�ǹ���k������u����;`�ǻ[�(5�c
���D�C���]ͣ$&��
k�8�v��3�u�ϰZ;h_������t{��W��	��H��Sb��q�ga0z?^��A�s8�w�03�ڎ2���ہ1�T�*���*kP��P�
�z�48��.ј���t��*aO��[��H��-�9X4����;aЭ���,�:*�,����T�>��bY�У�GYl�����&�%�ǰ����{c��XU�ږv�9;�9���ip!.�')�֛��s]c7����8g�QU��{7㙆.i�
4q.�P�4JBWV��| S��l����Ϥ�`\��M&�n���i��%MW�7�������>�3{#<��\]�c��M�@�/z}�OҢeg��A�1z�,6�57�V?��C����q�?6��6L�+��N�'VGA�oWj!��Z*HP��S	�$b�2��o|��s�DV=f�9 wBe���8� ��ۜ�í�4&%���~������y���#�>@qډ��Πǲ@XfU�u�ស����YOAR�'å.�11�>��L���0��H�q��U�C'h/���AN��OSO��������dxM����(!�q�I3���2�F����}��=54�[y���{�j�z��C(T���B��~����w��Wed�Ӫ���e"(YA
r�U�]@���xV����6�E��i݂�P���P��B�"�@��Gg`���� .hR��� �a��{�n�|�߂�z�ޑ����◲�;��l]0�=�T(8O���$�u|��J�� .�B��,�[����W*�
�}/ۘVPQ�fmf�8��(b�=�=��I�����\����s��F[P�# z���S6����p�B���������|����dN�x�v�݌eX��J̉�C3�ě79�GG��pm;��e"�����'��[�U8U6�o�;�t=#�}������ �Q�};g4T+N��c4O_��/�:ّD0����/�-��˯6��1<���d)#���[�ck�|����"FJ���
e�3�qͳf����+�VY�Ӆ%GH��g��`�
Q�9�X�ҹ��L&w�"�;�6�P�k�M���P"�{�߽ �0W�	zٝI�|Og?ݍ��h�1��F�>p�@O�5���V�;}:��0o&������){˞�"�.�{���bj�Xe��9/���1w?B�Ez@�NЉ
6^��:�w�!YR
�ߜTf�R�e�+sSVT|3���S�1ʺ�`�nzO_?`<��΃���m6��?�E�}�5�Oz}�{z�-uW���hImV�_]�샇ȝ��ll}O��E5�9�8�g(��G~~A����	�-�(�V)`p����g�JF��{�|�q��|�������� �YUP����yj�޹��4���^�=�u��{���ի�t�[*�^����� #��eru�p����ڞ��\�B?ZY&��e�〤ܧ�t��j�v���Z�$��_��Rq�WO��ߒ �*�����0��*E�K��!��WC{Q	��HO�-hlk]�5T�2���6���x��-��zl:KvkKü&}��c���D��s���C	��F�x��GU"C��P�M�t��8�Ҋ�N0oz���C:��7�?Aw��(qp �R*�8�
��=��{��:�r� ~���n��-�N�5��B	:N5Z�n�O�x���>����
��r�V/����б/�k_�G=N�`�"	��4,>��H��)���pg�K�ᲆ�����nx�@O~��>oί�_\#q�L>{|��kWA�����J>�䅘�V=���r�۵�+8���G��H����.�D;��cJ��i�&
S��>99���WA+��a�cn�ﾢe2��3�BX��&���Ҡ��L�ׯt8��w����� n��.��oh�=ǫӘ�F�$h0V-��+���������(�B��`qYgSh�}�<�����Bۭ%z"���bX=��������d�rL�%��);++fC��������PYM0�g���Ԛ+}����U=c7|IHH`��U-�wUȄGX�>=�8/qm���p��`�����&?U��[�oH?ϝ�h�Kx����uXP�ݛ��fu�f0���/%6��a&1 �C�ۆ��wmb����=��b�۳g�XAg_>h�dP�)W���e<�@�������܇G��S�s�����l���|��ys��f�%��mu [b�^�ŉ:~��i�?�ljk%bz�
j�,�֧�o	�:�֤�O���� 3a��Q��$\M�S$�D��[iXC��7><=����Y1ݭw�hi����Ʋ-ʷ*`�A��;�?xɶ�����8�3�7� K�B��+g�b�҅n6vK�!�<Py�Er��.Z�tg=�u��l�p��(cF479�ea�i��g�|B�<�����������I8<�B ����99�2��5��]�e��.�2��~���r^2BKӨ!��9��g�}|�8_����+]Q� ��9M��"�7���<Ck��t��FS3�j�ߔ������/$��30��x`����D
���<B�Z������V��Ʀ�{N�dC~�x���lgĄ���]P¯���u�E��Z�o�
�
�9��F{.�X��3V�1�׮d��v�eDr����1Ň�Pv�*����߽|T|u6E�_�gS�T�:��bz�(N������ɻ{S����7��-
�0f��y�l\-j��#wE�{�:�G+��;e��E �+Es>����_�䉗�ǿ(P�l	� �j�*�/=7`����o��z�R��S.:�r��Ux���_��`����%�����K	�)0W�w��W�g		GJ�}L��L�I��N� ��<��sf�� �[�R����qʅy�2e�劄F&��Om���eݮEQ���u�@����O���Q_�l�)
�g_����|MDv�to/�8�_�<�A��%8OM6���� i�k{y-��o���@��Z��n�?>;t�yFA4)���;㿛�5�~fa��ipgcj��:2�R?�B�(�Q ����������<=E��6=�B���)'�/ zSS_��e���oy�L6��A��3��Mn6���xD`Jny�'��Q�/g�d)��o���\��+����b�ws�y��H?`��AS.|n0#�NL<���bF��.��U��0��KY�Y�d����&�n���;2�!�r�����0[+4�*t�
+�W���\5�?� �c@+G	�e"�@z�XS}���1bڑ�7��<�-彺<t�9[S��$HyjQo�ɗ�.�x���K�.�>�@�0�����ou�0  �VlQplՙj=X-v.s12SW�Z��!9�!dj����o-@$�����A�=���ܞ���C����nM���p�m��Vg��/ˉ�_��Lp�����!R;Y#�ts�&� ,��m��JluT��AR�]�X�����3���/�	��ζ�P�3H��PeJ�uζ�ӧ�� k�,��	T�@zeL����%�B�Fg�[}"���)5���E���ȵd�� ��tY{�������MO�{(��)��H���C�f@�>���#�/�"�
�h?���"풠�5(,4;��b���Q���?�uI0�9LI�	����rGc��Z�$ ���%�E�S��bM��������=���>2���"45A�J�#J��Z6�\c+�Z�|��^��a6�7�9�Z��߀�zh�]��W�@�O�}����e`x��N�E�,���Hn`�:��.>�ɏm��UY�[7�.e��S&�U�a
l˘q�?b~�{���5�wiy�)��Z��'6���bbM;��^�?��m�{��C��o��K`{�t���$��q���'�o�y�E�Qgi�i���>�a�b7����5_EEf<>�Sлn�=��c�xmԠs�_��xn�Bg�����m��9��Tw����d�t�#����L���o3�(���SHTKds����s��o��n2�N(t4a���y�Rg���(�DAuOϦ��ԯ�l�J(]�@�zYII�T��O�f�"���^:���'H�� �����ҟ:O)W�%��0��J�+���/�"��ᩆ?y����U�(N�L���䤵��]�Ԁ��B�Ϋ�2�QU���N�n����
�CM1�nh�yʯ@LK*%:��w�J?+>8r8;]6��+̉���
],D�+~U�aץ��Tq'(}�2��sΗ��V�����E&�/%���HQ$0��3�2�0E����Z��߹�� Χ?>=���	G�� �^9����@A��T*���<�����[i��N}�ME��������ڋ�H�+����Yq9+�������Qg��7�rP/@B��WP� �K`"�D8��}��j2�'������cx�?G(s�%]��uF�m�߁��CPV�5(���F��4����y�w��Ґ���=�%i�^�Қ?��˨��aa�u��;#�����ө�6l��k_~b��o:���N��2��Kh�8;]!.��kW���<��&K����d��ol��Y������L��ZSb�'��F�2�h�����33)c�����|C��L
�o ]}V�q��M7l�����yk���o�yV�,M��Y�M�\X�4ppĭ;����]��� �m�!��*0����Q_G���a��E"��֕�}wm�����ė�f�X�oF����u�_g.��HLJ�P� 9n&��Omy��RJB�̳��Q����A���Sg{�C��#��A}Ǚ�>M��J(�e]��{�����;N��l�\c$�]��b��c�(��?դd��
��nݣ_?�1y{M)�F�^,��ʂ��K5~Ʀ�	�!���Q��$[+�E�e��x���*��n�	��T}iiJ-A����fg��o���/�N`>Gg�=���ӳ��g,Єfn�ZO~��o�}����? ���z�Зb�+N��Zx��`6ByIYR�?�p�� �h�P�4�/g�m�EJ%�.���<S03f�k�D�OG�q��򱎈���CS��/��xa�]���s"/�;<�<��6���fe�j��#1 �S�II�+�2�9A��z@�X��/yi��4j�p����NB�\��S�D��k��*� l[�߰���Ï`�e<ut�d��{g:<� ��UX;������'.[�I�K˿`���Vg'�ԖWQ�az�=�[\L���3��ou9�n�J��}`�_[vdH�7*���qw��k_�P����IM�{#��L���B�4ہ�˓NLe%^����W�-5������:vw�r�i�yA��.���{7�M�N���~�w�o�
p]������K��P_��|���6=�����s6?,����,ޚӰd����*-c���(rFZ���U���N�����ላP�)���0��!��rCX����1�(%G���g{D�����f�fF� ���F5rbH/Y}{��fcX��j(��x9�03�\��oL�?�g�ȭ��ѹ�ա�*���>����x�ԪE %�sfֲ��|c|�Է�&����HyӈN���>�ۖ㘺Øz��i�~�b"b[@p:3k�K+ ��JT�����wQ-2m�"���g�����9��g��F�G�����V<\�;�ʊ���H����Ր��'9-&\!���8�[�Ft�U0��D�}2�I�bc_�?�%w��7������%�W��!te�����Ý�`�}Tv��@�Kee"讞-�pn���F�q�Ag*��%���T��ѻ�%�z@�nq	%-����'r+�îO����8�X��Z44��7Xc`��ŉl��\��N�{ދ]�w2>1��wW �9����&&��Cx�!*����~�m.��=R `��=\�W*�j�}�c	��22����#&	���")�Fݵ7��� �0D+�������A(�)��"�������t���E���m�9�w,��$�:���#��M��i�y�4g�� �)�x���ra=� .\n���H�brr�]��:U���^.BMr�={��LD�'���֏��~��>���ںH�=�%^?C��U羺�J�J�4��X-o���&�-a�S^�qyG�r� o��U8(9ygz����t��A�<^�o+���~ �h� )�nV�����{z
WcҲI$@\>��&P�r�ZLlxF�w�30� Nr�E0@�Q��8/��3ߨ�_U�6�P}�ʊPO�'�c�$EEl[R�IG�Ԟ��\�G �	�M�0g~������tĒ��	3�4~�]��%T\�\[[BC�SQ�<� ]K��n�)/�
���5l�hT`m�?T�@ ��>�O����q���b'� ��Zv�#n�̌_F6E�H˪�~*x��߽a
�76|����� ���ٙ��+E��0��{==�w�J���B��6uc	o�;~��Y�蓰�ܜPK�nc=eO.8�n㮝��� �j�	�g��61q���S�Q�M޴q��Mx���*�W���. q���V���,��?����xy+�#Cԭ� R�3���ƹ�&'6c����a��Ҡz9َF��,-�����[��6������3u�Q~��Ri��:آL����a�3�D`�w���-���/�es�Os.F�YM�_��`�ژVJjjʮ�;�KX���U�X�y�EYVߨ��ӧ���`��~xϷ�"NGd��r��V;V��eώyf�,?�r�����jθgE�4��60h�ihX�˟Ů�<k��QSC%6P��ڴy����T{;�#�y���J�ӧm@�L�
�P%��h#GU���@C���^���(�+��x3��x F(�|g�D�&�;4�����Ol@�ژY, ���?����3{D�����+�!!F���Cz�m�L�8R�X3�ﱈ�_�'r�K�6N�q)<�efU༢�K��Oҙ P^�˜k����N��g� q�-��7of��Q^��{1���3����huqqs{r'R��T����5Wx��Bs�[8 J	��M������ǁ��Ύ�%���gϘ�n�L���VP~���W�+���U]�;�}=fqW��Q��Z��&���(-���-��"�#d�:[Բ�PR�J��l-?�VOF����t[�"��V�qY݀��D"'s��T۳A�>q}SS8� Gd�o���a�zS��c�D��NSS�Q-QSK��M54H����h(�e����햔:�QK��[�Y���.��Iʞ�rS��HK(-.ݨ���5� +��1eG%&����IK�{:��\]�+�?{uIw)X0��$�|Vt5/osK���+M��sdFq���sע� ��e9����d5��F霼��Rū#T��U����hb�ײӦ�aiU\\���s��C���q?ƿ8���1���-����)滛"=YY��2j��y��"��j�%ݜ.�3�'�4r��� ۝<DG++��gL��\]Ӑ�{��?�x�7�A� Ô��Êv�t�;;\H]��[�^_�������\�w7�ݽ;����I�y�($�8�ˠ��ǎ���Ϙ�q>�+���&�l�:u*W�ԁɅ)�XZ�Gӊ���hb�Y��zcs0�P���G";���8;�Vդ�[��Xpw���:���"]W�9����:a��yOC[Gf 0I�p��3�ᳳ."2ȧ�:Q@���x �'����H��+��&��1W���3L�'`�J�]*jmhx��7K\m���8��ZZ&����XYv�!�g��:�,]D�������C	�\��V��('�:zD��bz�l��j\VցD�DyR-6�jxT��zd�`��,�lm}��^dhh$�k?C�Smh����S���w����/7T�YE�r{*�? �a��:������i�.��z�N�LaF�P�Hg��?XGq����mxex:��%���33��x,�{u�<�R2]qeM�r��z����Q��E�`����"Q�V��4�/_�~��?���
����g�05��o=��ػ|p~ߺj�<�`L�����a_��z��Ƶ�f,��E<�%׿&����>�_$44(ܢ��1�T)��$�Dk4�X�.x$��Еb'|98��4�L'+��ϟ�%&�����$#������#� ϒC�ߟ�Խ(�0�s�r�h��W}�I�3�R{Ȯ��j���OK<b��	�'Z1�.�n�E3������!������|aAƊZ\xCOIT�p}UC?R������o��H����(T��#�m��}�T���i�W��1Pkt�"XMc��~���ʽE_{�*du��T؇��Fk7T׊1�ǖ�L�0}�ç�~��3��b�%{��!�,��yr�$�1����Su�u�U%��v����Y�o���}������*@�!<�jP��R�=���!�;!y���`F�o��նr�f�~=]��>�Y�c%�Q�bK��K�>���.��RD�t9�k�\��{�M4ΞF��<�H~�P鏉��h��k��Ϝ�z^���U���q:*Z\yچ�z�gzh{�C�[����޺�램��� ���i��y��**�����P�Oc�!��q)�{P}��>~��q�ܢ�U	�|��C����Đ&jB����w����.M�0�I|�9��b�[� [�gOk�/N8��p�v���`"�$D���҈�X�П[�Rƌ�ש #�?mja��]�j����@%]���߭�yP�g�3|�]+c�MA�A�ꡖ����iS����`��\�ę=�w�y��؏�*�T�u�Z�����U�ɑ���k��W�=����J��[���󈐀-���m�(�2�Z�x,�r���渹K
3����7�O�s�b�'-E�Yn(��|��_�ǵ�Ja��n��ǵH�i0��kt�JM�����
s����'��8�?[���k��v^��v������;������;������;�_������5	|�a�
���;��؏�[?�~l���E��ߏ���'�~l�����c��֏�[?�~l�����c��֏��/�.{,�����+�n���h�N\=�W�	׋1�1�
��xo&P�\���<TQ&Y�q"Ź/��ގMH��R�;iy��������˿~������N��O�Z�����1fj�]�4�-�+�k���L�a��I��]���n�B��������^�+���m���BߏS��������){]З�U�|�Y����7zz��꼨��Y��=�)�Yk��?}M�jk�a��S)B����s���������tA��*
}%���t�@õ�9�񋰽�,4):3B�*J`���B��e6�A��o6�o����k�.	��D���q}�������>���o��M����.n��+��8r�[�����.�yM���|�C�?<��}�qrq ��7��/�m
}�:n���̌��o�µ���T� C���IP�١\*4�ۥ��4�b���Ŧ�h�>��p�FA�����;ڧ�//]����tH.n����Q�O���E��[4:>�/�}ʇ�����@8��M�Pl��� �4�$������U�]�y�A߬p�ɑ����B�{JEK.�߾������LE	�7%lV7'����τKF�u�߰�y�;�d���z�ף㟣�V*q��/)��I��Z$��צ����C�B�����C���!�_@5���(W��(���v�Y���\��k��Y�i%�hx�r�?���e-V��S�8lv�\^t�W֣���|�.Q���#���@Ay�?v�e���VrBo�	�������YJ����Q~ڠz+Ep���;u%����;ڿI?��B�9q�M�+��4�O�(��ۂ�d�v71�g`�9H\Rcww��t����971��ndd$�C�o��7(+)q��⳱o�I��#��!VI��v%� ��1@����=�"**� d��e��"�ww=�+�]O��@�K�8��^�.P��f9tO�f�7�:W_,j�����C*����q����PY�}ee�%���;��u��e��OPS��0�L��6t�2�!�Ԋ�	�J�eqǑj�`��������M��	fbb�8)@P�p'��\�kI�G�D�8M]��4W�7�u-���� _[��g&*�nD�Z �С�Y��X��ᒀ��9o~$@K��S�FPj�7Pm��_�H��C��\X5�+�{�5�!ǵ1ƸlA`�����̲\TM��h�m�"�g ��`%��*����b��am)Z��ԑU��h;8�-类;��B��uG�T�J�`��1�a���v(��t|���V�'wwu%�(2QQ�	8x��M�]!��G��X�!��̃�ammmVV���Co~���  ��'Z���kӔp�ySllk?ӆ�?U�#᜸�?�`�M�---=�d���eg�/FO��srh�A'�?:�0=M�*��P�]�"� �ꈟ%09���T�R��M$w�|��&����C�$p��E�V�"�˰�K�vF�Z}O(V��ZN�е_ @z��J��<���~<�팘�~wR0d|G��ˍ�I���\�X�w��f`�SR�H�4�ae6iu� `���LNFX�p)B�q��8me�������ɷ}�`àOܭ�Oc����u�;ݎ^P�+{�1r�4����x��R�e=Dˮ��~@� R�;�ӑ�Km���ߎ�y�ǓQs�+�oBrr:2c���gԔ�$=�����-�.� *��/��P��Cm�8�����B���?c3����I��$��B���� T�6k
��Xv�@�P�^M�:m-.*�HPv��}�\Hs�A�ǀR��yH�� ;� ��"PR�R;:/�z�j�#��`o��	L�MR��?��p���S,����.F�r�p "�r�ɣc�b��b��N�-�'��GZ�w�h\T:�Z-�vy���G�V@E����)�wtv2�.1�j=�zn�)�/]����W�ĸ���v/{��2�̓71�����UU���j���l&EEyD�$�=B��� Q���#ge�+P2�1���=�	���Afi�8( �p��0P��%�Rڱt�g&���Ƶ�}TO���B郻��I�'��E8 ����mc8P�:7A��^��n~��ys�m�)Z�|R�yX��sH���K �� �')U:�<L��y��0��yj �C�2����b  K�{3)rEE��9!^8�r���k
gAX���J���f{ĕ_�컀�C}F����&��*�*�Y-�l�*�hY~mHNN>��Zh���#��azT��V`*ճS�h �E��������Ǭ�0Y��� y��׸pv@���U��tP��g:�JKcc#[F����815W]�CՏ��*F��h)����g�T�$��
���Gb�:v0�p`̗��!`�\>�.@����L���[���� <fa�<OL��֦X�q�[@�ٌ��1�Ud������Gd�����Ǘ�&
8n[����EnJ��{v�6���	ǌ2T���A��3ZUV��0>��z���<� .aąs��93:
A��:�D�޻�	�7T,��Mb�\\!vh�|��)��������J�j���R�`�TY�(Dl��\��@Ԋ"�첷V��P5
B ���,.,���1(����Md�fNr/���?��9sf��yfι7�l�w������..uW�Ӛ�Q/Q�����u
�4���yw����:��r&�OS�B�:K ZG�3	LC�c��(A%#�M�T�pG�a߻�fӰ�e{$�~[J$��эw34��'��\2�/�d�OԾޢ;]UXs�x7�j'��-�8a�!�w�}�V�ߕ���?e<;D^a�\汳��> ��j��3��O��`)��}�١�|9
j`��N��)���7��9@�f���`^yY����WhlM�&P��'C�jzw�H}9����w���9(�Jm�#>��&�߹��G�-	�-n�6֖���4=Id8��f�~��c� �u�x�<sΉ<mA�:K��[?ɉV������i�R,��5&���$�DSe�YIKe��1��`��u0�qǿÔ��2�!�q~u1����n�A�xa]�%�Yi���D(3uJ(���_��16�i^,�6��v!8�'�el��$?�)�QHXN"U���DW�#��Í(S0��[wz�����ˣE��d�4��Ӣ
=���O�}R��*�}q��I�o��(T���zZ��)�7���95������w�/ 
||�c�k�J�3���b3���p������R�c�w˥�͡��wi��T�cPo�|���`�zT��vH����x�wO.��n��2�ǒ������\qy���3�W!�m� �Rh����@�]~2eTT����0_*5���nB��[˲;��(p���~� ��c�_W �E*��E��2e�W���ڰ�
)��z�ѥ��̢i����
K&�<���v���nkg�%���\�%~i���B�&&��A�y�D��TŹ��սc�"CD��[�0
B�)O��o*�}U�ݺ������2)4*J��x,&L�qGam��/8�Z�6D�oPk�=��!���<y�$(f� f*z+D�����HR.g\����m� ��<�,0hEzMލ�ք�d��x�rf��4.Z�F~�K�+��H׼�81��]a�oE�v��G6����'L����e�T��>���N&�i�5����6*���h�y��w��#�^����.q6E�Zq�_ډY�݊�y����5�&[�����`-���_Q���k���E��]�Zρj��]��={��5$�S6�d9�o8�ϝ�s��z�m�?��pn%�ХH3뚛�k�<=,��>��R�c�����
=?��DD�{�מ���2p����)��@=^�y-��>ҁ��{��3(�����
[�M��y/�K��j�;P@�"������Ԯ�\�Ө^ZX5�t��"7���V�e�ye�l���?*T`�l�D�3���.R�� '�.T�3������_PK�C�{�Z5�{�H��gKK�W�P=�/�۸�8^������%zz��I�Ĩ��]�($_���8�Z�L�$��c���J����T�[ePA�W�-n����i���m�YMt��I_�@�h荨b��҇p~�ܨS��䘥�U6l����DS��!//��I��d�T�*�z�Qcwp�p'm,���-�I	�5�F�k;���v�Ռ�u�?�ZRS6t@��+��%}K̻��3�+"㙪�S���Kz� uv����A�l2�q�בV��<��dk��z9L�Z�
'�n�R���b�4�w� 1)��rp����gz=�?IzO�f�]o޼9XS]=C�`��=���C�1��B1M���׹��5\���'_w�b]o���I~5j�t׫��P��u�\ۼM��(USv�p��p��P:���{E�w�׉�r,�78<�y���i
����Q�\��&��+��`�IB�u�hx+���_�����eb9���'�QķG��wqr?cD��Hz>%:5�`�0���ҝ{�t}U�D~��7����	�gɦf*ԸK��Hw� ������_�>gK���^3a�u3v�,p�h'�x��J�H��aN���s���������lIp����)֥�pmF�E�����$4_Y�Xߒ���Ιk�Ԗ^?�e��`5[m�$��)ƊL�"�Ҁ�����89�e�y���X`kY
_>s�����'�Η�c��}6�}b� iU"�Rm¥�Ӈ7�Z��N��}�.ni�E.����[�,;�ߍ��]��<�c9�!�Y)��8�Y����$�h������H��K�4}iU�Y��@�tॏ��Y�9/�8l�x�m2�]���Q'0��V��?�1μ�>�A�;�dȰ,��H�i�ĸ�E��^l��
d����o=^��-�x��	n�O"�������M�F�6v籃�mR����(����!�W�T-f�3㵼��bK����))����E��%دcc	Z<uh5��"��\��s�=	<.��J�������C��į�Q�L���c�!���B��jL�w�<L������X�$��5+It*�����'��LU��� �P�4�P��T�"��������q��I��h�8ހ��c�C?Ț8P�
�$b�2���<�V��S:8z�'�u�H�l�_X�o_�4���?Y���{��s��7�gXֿ�b���{YE���߮NO[Z}��__��u��k�������W�t��/�}~�r=�.�L�c�qo+?�*è�Vm�ќ"���Qmc���_+@V���]O�
7��}���i��ɓ'�$�i�:EfO�BG�y5'�[���wg�tΘ8~�b�=.ەi�~X�g
�K�a<��d���p����P��WۮA��3���jhd[�#t��-;������{�"��[_<��\~��օ*eKa>�$�$"�G�)NH(8<?M�H>����4�./��H=���7���t�yc�#!hU�i�����[�N4?�w��؅n'zӷ��v�-;Ў�AP�w=7�KGy�)�����x����H.WhAƪ�(~����F	b�ɅB��O�#J^Ң�$���P��A�nQ�-�����"��ϧ۴���~���7�\S�Qk���ؒ��F[H�O�[�`w��fO��zG{ޥa�)�l|��Q�l5�竅D4�"
�{��ʤ��?p��W�,Y�`�<��1����\nQc�!ˍ�z57��-Mt�_O|w��rc�Н����"�kɳ8��������(T�⤶ƢQ?O�٤1[�}1��9b������L�|����������}~V���Jr��+[����-Q�J�vg%:i�#1cTQw1F����0��� gWȒ�---}iJB�_�mHN6fv>���gXT�co�=٩BgM�=�Bg������Z��l�AvM�y�ۤVG��p�� 2��w�L)'�b!q��J9�� /�]�h �y��
�z˥�ÞQg�ImO�Ԭ*QC��}:O�(A�+0��������M�J�f.�!L����O�0�ߝ�ȑ����*<����AuuujP�9X�^ÞQ�Gb=���h4����>cSJoa�S�2���B�z˪"�������lkW���6(�V��0�w�z�č|�ԙ�o�O':��)b6���8�F���-8L$��6ZV��SF��@Ss؇;d�>|�pgHȈ^�*��3��*���ǎ��Jf�������J���s">��(l�Bh��_�t���C��)$x�Q/�^7٤��m{�YfW����:v�<��==B؈���|�Z��|�L��,-3�B�p]DP.*�kw;���s �MzxyQ7�Т�Q(�F^�d�����k&�=�e���\[�����k���]ޕP��N��W�������G�[����j��A���+E��|���~X�@��8���L7�����ۥ0b�
��w����"Cm�w7T�I|~I��gݻ�Oij�Dyo�E��?�5�)�h>��kd2�������i�iɻ�H�xy�����s��
GmqQ�o@ na��� �L���_��u\xO��ΓJ,���y�u_����5f:��5nٝ�b��'!B�Pa4Al[CA [�s�l��GfĮR>j��(�0S�]͊E��ڥ >1-
�יe
�?5�w�fGp�ߨgv�It�%�,Up�����B#-�<t��s��?>o�w2g�H��82�/��v�^�E�Hff��$uá�D!O�R
٨�#���dN�	�yCh���a�}����F��J�1�F���y��Z�p��I�����W��[���۲��݇��B2�<#P�w���O���ų^!�v5F	��)�1���ʸĜ��ڀ��;�Mir�Z<1����������s��c����ξ��J���<(z�B��)M�1d�k��u��������I�tY��޼��?��#�>&�`^��"�����+dwhF��{�5(�-���P��{ o�II�ƶb� n�N�-�R7�����N�vVjʶ3P��L�(�Rw7B�@��G,�R��J��T�vR^ug���ѣ� ٜ��Go�Ȣ�޻w�Y�;��MwJ��4�b���No-O�wk�S�G�9����9�L�:/
s!���w�.�~Se�hNg~�)>�ȂL|�Ν;��z�6
�)��%��f5OA�S'7>��QFB�E���4.��aN�?q��?7��tM=� ����V/�	z��"~n~Zk
E0���@��R��F�w(Jk�����J�MP������)%S���i_�Oi#�`��	�2<��n��^���0ϙK_î/��zK�WG�2)
��C�ū#oƐ2G���3�����������\!�+A��S�%'��L).�ް�s[��nS:2<8:[�3�Lff �0�ܲ�����F�w83�u ܘ�%����Bn��u���Nl�
6Q*�I�n�r�װ��ԝ^�P��bD�R��?��s����� �`��@8|�[���(�LE֯3CGG��sFW��8��fܺ�Z1��}�@]� bX���G�{	s����2����K�9�(��F���{z��$x9�A�6�T��+n^�}���g4��9�k���Z	6�:���DR����{�i�&�,�Ǯ������|f�)�������J��k���v������hcJ/� ����:@ �qM6��" (Fg�X�{x=�ŏX�v9��
�b?S��� �L���H6�a2A@�,�&�b#��
)kZ���!r:�9���l^���j����H�#�Ϗ��n*�P�u�'��J&gj�������^	[C]��X ��|��<U&����D\s6���~M�dB���#�}ɑ%eն���4�6%Z��0џ)MR�?/��[E�*��O@/�k|�%��s)LW&)�Zka�ZY��j(�] �;qK�?G�l�k�!cѫ_���5���<�q5�)s���d�\��=��-�1��]MԼ��Q��\}�5x����P�&�υ�VO|�_N.��_'1�'?���X��iS~Dx�tt�b>� ����Eɕ-C��1JO}ww���aP�5Bé.]��z��l;;b��n`샱�7�֧��G=#�����A�Uٙ�oĝ��G�'&֢L|����Os��*�W��v[�:S[?���N݁����v54\�)T��ׄ)�������BC�@�����b�0����=SA��h/D��Ľ��Ə+�M�i���9����[&v��}x�#ۈ�ϙ/4�(hx!� GK�^�,��m��0�.��OtvvN�b�/�8%����]��,Gi������@_^�v"��555�j�N&%K�%_�O�$j����qI�R۞��Vc��d.��R�;(��i&%	�o���q��IwB43�Y-��MgFa	�g����N�9�	���$�a��
�F6sU�=�SZ�Ty�=���<�p�I~i�o{�n~"��P"JKk�t�`�EI�C����Z?��� _���?F����@F|��-��"�\'��%m����9��ߺu+��0��oi
�6B��_M�I $������3�~
A|rg�7mU�1~�����0\��$	�n�on��s���7 �����f�
ןFk�0��RB�pB-�٘āOıwRO	��P��%�%Vp���ɆҨ��ɅR��Br�^K�Fs���-�w׎�wS�;��-���4�73��)n�LOq�KS|�mo��#��"��%$aL�1>/J��k�����z䓡[G'����y���3�/����h���_-n�ĴM�9�52"�+�/���e�i�0G}[Pw���5iiD5v�(����p�h;G�4�o��rVH^Ւ�$X𲡸4!9��S�����i?�J>�`%�x�L\�:u���qS-Ε���m����>l�����Z�Qw2�����Y�a�"}��2Hm)��n_��If�C>m|-N @�! ��Yi�1o�[3)'���6�Ό���H�풉C��bn��(�S�l�6��ajL?�dS���s)9�m|�Mu�|��w�K;pQ,'I�=�ԩ!c܀���x���+[b�힦E k�@��Χ*�"�N�����3�� ls�dq~�o�U"�v<���z����e��L[u)��
�4骵�:�;sq�VNS���ýGz�e`��uF+;R��?inn����÷�l��M���JNA�i��Q����?��>5�y	?0Ց9,5���լc��fz���WEE�qS]����:�+��Bф��&YB��q��PU{�{�^o&k/���.�l	�͊��y���\�5#�$#h���a�?B���'��&�����Cjb���s
��7�=䌨�A"
 B�E[�Rq���l�N(�Ĕ�B�dh���S/<�Gaů��v�&�&p�t��"��N����fH/��	�R��g��<c��1��0DކA�̉��c�|�8����Y;8�ػw�I�w��Wf���5P!b�f�۽�L�V���B>o�O �lV��.�{kJUn�SL��>�C(8�@K�M����K枕h��-C���XE褛?�9k--[������b'��L YO����|K�р�C;%��$���$`�v5嚸z8u�A�Mm��{���=�nu�'�D�&%>`���J�����ԏ�;*��|Α�,6�$H��S4��{4iۤV[���	pxlY����|�xj�K���+��3ձ�W|�x����d+��r�gX��ˆ��a���/l�F���|�B���#�P�Bv}�p�����-O���[Ba�*;��0`��=���7�ŷRU�z�z��I��s
�W~:6yv��[0kͣr[��6�-9"o�0�z���:��G#���T[B�*��#�SZ>Y����s���K�b&�춃�Ozc�C?��N�h�pܫ��0rēA��a���6~ˌ�r�Ġ�;��GIc�4��Rq$��#B	z�K�J�^����
�d^�d��ifl��d�L=��tBXۨ����ͭҁ��Q	q� �J�u�]�B�kN����,rP��[�����I�O�h���M��`��/ ^>���֒0=H�bQ*p�]�-x�f�,�+�®F����dj�D��3�v������π�+��Y�=�{�����D�3=�5��B&�\Q�	�>��$ޮd�O�J2�b��iK�o�,�N��e�}�W�)7W���g����)��׵���kB�4f�x���.���$'_��Ѳ�^�{um�y}�:�J���F�P=hM/*�CS�S�|}��1,��+��m�"Ɂl�×�@�mL1@[&xI�I:O��n{zE�Y}C]�9��j�������li�7/؈�?a��[��=X��G�)t�*����#$J>�"��/هz�C�����.y���7�=]�3�ض�\i�W߫B:Ŷ� 5��8�oyb�l�7T6YY�[#��_Lɲ�wa���1#��~�z4��#k�/�B�%�Λ������P@�`:��sێ���9�U�h-��
�f*��s���PX�Z?��P����ɌMh��$�K.�����'��bz�zrO0/ �]�vͮ�g8H���b-�#h�˩�P<�dسK7w/���J���U��!���+kb?���\�$"h�h
)�.{��9_�^8��K����9w�x}�����O���̓�-�P�7��}Y6��V�6��7�~��w�p��`�Q�<9��IĤ��$�PW~��ݯ
�g�G�>���H�ܑ�hg
~�+�k��2�&���[�6��_a�ap��S[':n|>�M�-oFۙ��"Uf	j�WB�8�cJ�L����kZ3��1��A2�2�s�W� �� 6�z�fiE�͉��e��,�#_a����Ȏh4�N����ѣ��e�T���%�=�0�ҕzK�4,V��N���)�b+��D�W>^�ũ	ƪ����xH��	
n,���xw&Q��l�B�F#��^���-P�O��oM��.�+�ܕi�.R�I؃�t�;�%�$Bu�����YR�^�2�О���@wz���!��<{�<v��t������.n
��G
��^r��cK�ÅE0-�	����Q��Q���i_vm�\��0z<�����9��&`�{Xe/SSSup�u��XA�%�ʕ.{4��e�)���eo�ī2���{�ؾ�e=D���)�	M�zܡl�[U�.ǀ	^=�T�|� �eS
�s�@��	�1�N��ìq�:��-Abc�z#�jv�������y~E;!�_Dl�S'a__��WS]=U���\������hkkc�Ǒ����d�Fë�]�H�+��>|X�Qei�0�����M�Q #S,�m�YV�n�,��Fq�[�O�5ڃ-�k��zȩ���y���^��:Z[@��wߔ/_�ͫ��O�շQ�c�ՓwI�yC�ȼB>#�w�<�传�w��)j�ͻ-����\���u��B���������P��W���R��F���?��7Ae�h�����%}p�ZM�Pi�Sւa���k8, ��z��*K���Hl�-1F����Ta������*���-`�y�M�x���vÅ����n�\y�'�ƿ�fa?^�~����]=��d*���rb�k&8�W2܁>gsK�L�y(&ѩ0��6����x�O^���d�t@�s<���1�5BuY��E�q)�k��=d�z�F(0�:
�I���@'?逦��9qѣW����y��m�+�H��)�,f�6	fv�S�Q��ᐢ�G���;�r���[4(^����I��9N�3|���f�1���+�1^l��[�W_U����vZ��-.NW�{%Wzi-k��+����J�&W�������w�)}{c���7_ٝ]�W��{��O|��-��EM����}�hZ[�Z�� ��s����t�\.׮�[2ͤ��s�{kϑ�iji��`�\B��#��o^Q�W�/W��)��y�!�(��H�F�Pb��MK7g/�	�/�a�pϓ'Oҁ�����ȣ!r��h����;{P}���ȘD��s����p���	}�;SzX�M6)n���É�NY$0�Rm�b�w�K��U.�.�����e���?c�|P͔�Xwi``������e�
bŃ��-�Z����@)�Ng�2���:����x"f���h�$�Ň(�k���ů�n�['�����Ǐ��kɄ�+T3�&A�>'�"}�`�̾�q�
3��2J9�s�]���cW4O�O�n��_��;��e"�gZw%i���Dۈ����I�j��"�Gݻܐ�esYD�K��| R�%�vQ�����Oâ���l��}7��?��G��O�v"� ���2�HF���ħnj��r�Dۇ�Qq�8�b����O3���;���԰%���,����LOK3��e���a����m�ήtw�qLF��2����C^O2)9H��y:>�p�L��dq;Հ��,�K��ˏ
�m�%!�+CE���)�\l���7�K�d���%IhMJ��2��$nn��+/�t�nS�D�	��}��>*�VBIfWc�m��B�y�l�}��~�ŒU��V�/V3�S�-���� F,'��+z�KK&F�B�m�<R�dxܺ'��(��"lD�o�*�qb|���
���hk��0�]��Y��`K��ml�#��Oe�L ��Ni� 2��/���ܼ��ſS�L���Ȇ��
���6�5�N�!kS������r[�*Q'�t���Z{?�5��R�{Xx�I~n>��gI�U���s�2t+�q�J�}n��Lt%F�P迣�1t����-+%����<�y��$x��0i���GK��a�l�_���WX�S�Mg[�`���i�]nJ�Y+ Ch%gѻ�D���C�&n��m��^.7������G�Oa`�[H�χ��vNR7��So�g�����*�l�ӣu��q/�̸� #�Y��{� �ߡ�7��ٴ��,�Ƒ�
gt�o@w�
&,Iu1�w���l��nZ�2_��A�"�!�|�:|>�FZ�IO��Z�~�?N��`�D�5֎�9�k1[��(*�>��/u��z�@+����Q���n}�h���Vd/ɢ�un�S�+����]E�q��k��a�k����bE-c�>L�:���t5;�:���^�w��<O�+�% ��Vd�c��7#}Q���R�Q5���o�BI�s�͔�!�v��ck"�1�-�v�q̬lɟ)���U��)�8�t���Üv�.��	~���s�4�[(����Ȳ;��t`DV֤�NMN1`�Og� gvF)=5UmW��)�՘��v����}w�Kj�
�x�tt<�r���Vt��	�Tb�&)su�<���D{���K�F0�"/)9�|^�	��2�f"��b��K�y�F��~|�~Qs��3tJw�z2�1E"Ga�V�/:J��PJd!�'��#E,��hG��!�~�Q�;������ %=8��\�%����*��VI�WVV��e�b*&	���շzJ�qK���Gijj.?�@�M��UM�mj�T\�d�[6�@���u3��"B�ڤ��)))I�J���%�Pe����=��:�g:�%x��w�����
�������ȓ(#���p���%
/5V����B�ק�R<y�^:
x�^�^���I�m�=[F]���֚{�3�	h��Sj
�.�*����)�0�XZB�;:��W��;���FԞj��6Z�6�|�}A�É��e��>�a�ǁ�����c�y�6�r{�n�ڥ-�)MR�E�C7��bF렶�𒪓�No�7^P��_�9#�!�~������Os}Z�k��v�� ����_�񸮮�!đ(/�o��Rw���WD�\G �����(�{�����[f�~/��^i�Mu-MMW���朲޲j��c�)�i� ���N>/����m��U��f�1�'�$j�K�4q�*c��`��-{�9I�I��ʀ R��O�}*�����KU�լ�lY���D�~OX�㟢�x�,--���s���~�U�kA��L�7C
��c{m�i~�w��Cn!)r	�8��gϞe��>����b9��r�,�Zc�Q�̶�/�Z�������﬑XV	3Y;��ބ\`�)�iRRC,x��S�w�1If�P Ly�3| ����@n/������xe���)�>���ݭ�]Ky��ƺ�ӧ�Y vz�W���
	9A�P#�A�Ѓ9@��{h���-tڱ��}�,����&n�ٚ�zrp1�����z_Z�U%R����I�ۏI<����]���LN�eItU�1;����ӧ7/@���%�I�}Nh&����hIͰ�*���?�5O\`h;�	�6����>��C���_p����H����*=���Oڢ�=\h5�x��	�?�*Lw�J���A����"�ҳ��һ��W�T�tu��s��/�<�����7�dK��d^����x��{�t�$�^J)Z��"2eK���Iyâv���T��G�����w�"��
ɥp�r DiG%[x���	��O�~*�％��qhѐ�~�wL#I&6�I��D��H�֯�Z��^����+>��wEid��̖���u��o�V_I�Ç�u-��'��.x�J\�?$3m$'�c#��W ����=�'3����99����t���PM�s�|�l$��͆-il�0�r/̖�ʲ*��yVs7"��^��4����YjH���8 ��!KEa�P�g>/��oP/�QeQ��+�}*���k#兑�,�����[�v3�m��r�����z��t���ׯ-�΢_�=�)�*9�>ګA�y��U����2���R�S�̄R�6�Bq��/q�94�ï�,�����2�ZEC�1,�ܧ�*�RgSJ�EaN!�W9�=i_�H@��tG�ֻ%Le����J�`o?��h9QJ�`N	�i^ҝ�J�s'�x��63���>v�סd����GF���'KD!EN1��:A�9e�e,-X�vr'��`�yqwh���N��tzN��v��1G�+Q'6H�Z��\ûh�ik}]�������*�Ϋ�o�B�v�B��sꀗ%L��I�\h�*���ak��Xc� J-̮�dM@�*�}��N�^e|�d�Z-,,d�_�Η,�0��:Ρ�	u����T�U�,�ws\���Ȩ���5>�D�Ә&D%ǒ(Y���dVٵs���wĹ���)
-"ϓ��Y	&�jw��@�>��Py��%$��]�~ɕ-A��݌�ɆHo�����.ج�!�zD�����Ѕ����{}p�y��ڝX��N7�����5����<�/٩G�M��dD�K�������/�|a=x�z>,A��l����g2י���ٳb��-��lTH���SKK�#�J�frV��\[H�D��MU�!i��nj��>[>�LM��Ԇ*�Ϲ*[��|�ߊ����{�����0_J��/����T[ufƆy�� \���3L`G�a�o��)Yr�oPt�`��=�r,0��ݳX��%g0.8>�}(�����n���z9/99M(L2)!��rU}yP��+�.i3f%'xI�T@�ܷ�0xP:K9L��9���ٵ�2�S��䔴rGw���*�cդiH.�>���~�.* ��H�FtI�����p�KLyN2p>'t�C�tl��j����z���NU��ʽk���G:�y�ƭd�B��K�C�� +}e�Q~FqbL\�]J��Y=�)���uq��9���4���eW=QDV2��jM۬-���cc���I�3�5	C���Y��S����ROi�Ye���ߌD�1���H��}"u�8���<�L�*)'3��(������ u��������ڎ�`�r��kkk��� �J�~�Q�qdA�x-�ɰ��:��n!MT܁c���������wB}�k�)Bs"�͂���^����ID�$Ok\�l^R�&;@���Ν5`�	�RR/����ͫ�F@Ѥ)��Iy�~e��*��%���3lQ�ѴvW�''�g57c{��)�7���83q-�l0�Q��F3�ڇ����Oi��p婴����swϴ���d�>/��Z��ݘ��ԡ#�1/�r`W��:2�:��ws�-�����Ɇ��X����[�D�Z��*�0����y�Gp�+�4��$=�)���~�����$B�3�eH�B������0Ԝ�M��B��k2�$�g�^fW!�Q�	>S��m���W�W� ��$>������>hb(O0�T%��%��=�3�����Ɛ�hC]Yh`�������4�)��|���m��Ii����E���yk��U���Y��H���=<ğ������yb��B�B�y�-�B�ZF��O~V��Q������*!'�w�} Q��	ޑ�1w��jFX3ԙ�İ�eG>��χ����C>ݝ	�E7�zDT�u��3[�H�b>R�
��1w�¶?Z�n���#��C��v���N^#���X�pA����:{�厴��6.IB��$:����<�L�Z6�'��i\B�K�JB]�,�jL�8|N56�@A���Ax����=��s݇��cS���k;��6YY��Z ��������0-Z�og��Cq7��k�Uq(�W�nT2f���۽���̮,����6�m؝�F�r�=�T���aNJlݟ�`H5��*�s�y��h(�F�Q���PP@����C?��MOi�۾����u���f�c[Yf.�5�A������G��<�~��߹��(��Ogs�sds555��Si4����M��i"��6)M��(����? a��0�lo����vt����|`6-�R����*TT��,h��C�v@��1�Iku&w�|�ip((�&��)t0��$�k�%���la�k�Î��K�2�W{�)&R=|e.xρc�e#�===��(k��u��o^(������tP����g||�?�kqT�}ܒ��m��Vp�����TQ�T_''�+g5�[�3Y�{����E�_�*cRr�&����%�r�ȧւ�I�p:���\��x?��Ǘ���u��yG��)~�牀y��<z,7��]W�����5"}|W���ں�-��*��[8�����5�3¿�;A1j<�ѱ��E����i>��k�tP�!�ʀ�.���Ӷ����������	M�
1ëX_��ЗDlkC�V�rZkQ����D���'���ebL_����7_oY5��܆���4��4<���� �Y��s:���]�K������k��o�U�Yv4B��ni��յ�1ޯs9�)%31<6b��&�.A�}�%i4����W�2M�NF��P��台�X�l�jV%<`�Ѡ?���<��s�Zn���������~�� ]�{1��hZjj�Ld:�٢��-!�����������|��BE2����3Sa:�!�z�z8�³5�E,��+l:���#H=:�IkzVe�福��x
���$Q�r|55�;��
�Hm�x�q���K��k̝�?GL�f��>w)?��95c٢E�9-�^6/BM}���e��w�Io��~~>��\M���KC\�٧n��8�=����e#������"��y�17 ?�_�~���5{y0p�'�4��q4$P�8�T�ꄃ�z�S�>���_C�p�t���t�UL�M<�3�Y�����.7�sFX_��liiI:1vj�P�`i�wb�1��<��kZ��C�w�eU��R|�Ӈnc�<A7�%>y�)��n�XOybH�����;+�j ��!��VA�jYN�����'>�\�s����Pt�c�6Ӣ�Xȷ��w{�\(�/�c\;(c������ҒٕZ,��;�[�0��G�%��D����OvgگǗw��*�~�)��p�_��[�C��*@&4��ݧ�A'�sbbb����k�ل�ߣ�`��i�.BhD|��h���#,�Ǝp�ִxO277_>�e��EY�#kO�������M��u�bSB&6�'#���R���TIg,[�Ty��ah|g?�2��HGG|�_�	���R|������ii�Ȳu8��昁ǂ��d5�8a/��!��8vj\�f�(l\mB/\��D�pb h��}�FwH�0��i���I������,�i�6!'�=_6dj^9��>D��YNn��<IO�P�@�d�ڬv쀎P3f��w�(p��jw��V���� �GֶۓN�8��Z��
�N�;��sxJ��'k%���C!k
�iI<�ÿ8��
8�n�R��ͫ��w���&%����%�˿7A�Pv�14�����/�{����IY�m[��U:�z�����7���w1Wk�¬�*,v�W�ε́g�.T8F}}�3%�~�u�p�x�������C���Z�̼��;�����㠾�Gy�95����/;��[��������~�e�n]@��4�j�������/�yٵ����y��w�ZeK�6��UP�?t�/޾;�MD"m�0'Z�~�e����T}����.�Y�Ź`kF)Xm��m��i]��+&q@��9�e'h+������u���RO�0��u��.W,`�^4z7fgg�U��U�h�=���7>�	�`%>�d�ȝ��3Fq3�M��Í��N��6�1�*������hS��-�;=.B��;�ᒖ���{��~�Ȱ���3��Uf�q�ƫ�� ���`�4%	���]����3)QB9U3�����E��U�����/��̄2�	K�k^�����J�^v��4v-`�h�U*��^i���������ސ��O�mS�7i���Zң2�!�ʀ�>�h6��XD����6��a=�m[�M��+��o�{��jq6�d�͓~���A�f�k���\Xi�3p�!����ͻ#lZ;w�nu_?y��4G��t��X���F��3�.=۟}���V�����������*��*S_%�N#�}�����b�椇�!b�:>X$�]n��BՋ]���O��j��Q�K��c�M�zt0�T�l$Ҧ5��u�[���6f���G���ܒg�yq~SOK����.J�����z�P�F�rS��G_Jtj���`�d�����=@�0��wcn�8����`�����������?�e������%��x�J�q}�����\�2���k�x5�����=zT	�vqfu:*e0���U�Ɛ�������$�V�msO���	'q��1�L�Y��q��98�σ�jD����.�\�>m]�N(�+JF� �ռ�|�&5�w�ɘ��$O $Xp�tA��]�9�y	�(}7��t���eqkC٬B�e��i;��;�f����O���'pDy���=�ڷz{{�U�8�1+�· |d�`Ct
;�OdV7��"D���\z��Q�"ufgq��8�;�sW����{%��;AxYz�n�D�hl'��lݠ|~vC�U�7*�N�]��a�>�	***�?;����^���8�C�|���q���� zm���D�pH�\ߣ���.u�Cv諎��`ȓ�ޏ!3�޸�C׼��@��^oe��W1��(�,�ruu���ه./{u�$rF�H�(��A�p�?2�ќa�xJ��$"D�X\��S�|E䩈�w��[���骯rA����}��T����	c���.g5'\���ާ��
MTO7���G��S{�1����<|�O�l����
Kޫ�k�%QWQ��?������z��6_���6Z��f����^Wm�.��ϸ$�0�W�W0�L��,����2��U��M7 ���0���ᶝ���(������#�~c���w#��N-��t�B)��>zl��ߦdV+|�	 �i,�f<8���16���in�4@�ر�o�x?�95���-�	�f��9F�o������r�����94�O����<Y��x���O���-2�s�DdeR�n~j3����3�gc������4�䬉z��I�Y�ٍ���+ �TU&�s�H�=�L�\k��C-�u	(ƻ�g׬vB֮�>����O^UrH����ga;����G!��5K�S���Ts\����ɘ�\:j|>{U	�����o��i���'�]7p�X����x1��}��DoFd6>�"�:��Ym��c��gli=�dA7zbSp�~b�@�?�[����#��A#l��;�c�)
����xP��7����������z�֟#��h��	�:8�zn�����D� зy1�{�ٯp#g,��G�ؙ5����>���,��������ɘq����5�\n���s?K�V����$�1�7�YѰ�	x��`Z���s`\~�J��
~��e��_<ϊ�P�pD��L��^���7:�}6�Ψ�ǐ2\koCX�G��3��q�)��<H�S�F�ӈ"�0�K���K�
g�F~�k��~AO��?�Ҍ��3	q�Ol�I�9&�E��zzf,�1ow������Tvz���|�Ljc_�ZQ�Uy��1B�y ��Ŗ����/�G�u�� -�<�ƿ���
�h�$hث�G�Z�p$��{F���f߂�۪���-��?�G �+[R4�ŀ�u�vw���
Cz��J����Z�|M�����6sA�����1��c8�~�ͬv�$��,�d�1�:�N��Ł�݉՟� ��Km�n�<���  �MA�jL(��:�kٯ3�`Q�}�$豵U�t0�rf!��g]��hn�]���e�^^�k0Fi��}�km|jf�23ҟ�R���FC=��3�V-C�+R"2@�� b�Y�����j��]}8n=����ZSX�k��[�� <�-^�������C�;�7��hGe������2t4vJ�{�l͂�-E�:%���ڬ�˙��� �܋�˔�}J��.����?u�do�������K�@9g�����c[
wuqY��Đ�y~}�������p��Q�;��g�%��w2+>�����ID����&m�?��\q������\2�?�e?����ask�����7}�q|���wà��N��C�l��683����C�cf��R;�p��~�
%ج��+*b*�Иd&[���{�p������|ļ��`�TYc�}����/[veuM���`?��K��s�7�﷏�.8��ӳ!"ݣ�C�ZV�Ǔ�R5P�߯�C��׎��rvn���}9�.��xJ�ec��
�֔�ŀ�]�n��P
��ql�Ū�� /w#^%6)h߅���fm�;+�,�� 1c죌ǻ�Cٯ�A&����g?����@��6_��v�7��vt.���k�y-���L$���%	Z�;�4�/=�(=���^�j:S�I\phX�}%���%��5��r�~��� PK   ���X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   ��X�A�x�L  �M  /   images/a6fbdf8e-bd4c-468a-8a96-d55269d19ee2.png��c�.L�&|�m۶mϜ�m��m�6�ض}��ض���c���ɷ?:��tR����H%)X\X  � #-��4 @�!��u}�b�'`��]  X��3@�]Ӊ�[�q��rU�m��a�l���`�v�u15v4g��l�}͏ �Ɉ���ɹ�
�S_�.O��ZO�,�Z��N$%��U��)�/̟�z}�	 U��B�AKJS���5�6�z�O�lzS�5ٚ�=���\�:NrN��R^����VV$��eP�̵����샿��Oj��2d"�^4-��J��(<���LLL�����7/�����>��=[#��]
��;v�};���3nZ�z�?r��Z\,���V�����s:NET�n*~����U����W,X��B#�z����ͼ��+V���
����^ouM�<�h�����/�.���Mu���a
��G"�u[o�I~u�=yS�k]7ce8�|��)�q�xZ��{����-��<b�>a`���� 001e}}}-%g2��%+C�@��Qw�yq>����	�� *���͒Mk{�u6Z����ܕ���R�1��>�n͑�U�#�S��^�ԯk-��xs5Y3�38�7Lsj���\ߎҁ�u�Y�*��h�$�	�B �·I*��ky��]ڍ�_�r�YcMo��������k��]����n1|ب ɓ!��:�@]�7��9u�
�:7�s;
GQȥ�䌥 ��#�憙~`�� �(U�o)3�Q�*wN����:��Or}��քTc��_\@X�gT���{��:/3�ɍ�ID�H�~<_B�BŁ0�\���k��l#��,�k.�1���&C��� ��b���N�r��F���߬����8=s0n�+|�}v�ҫ�8�	�@�T)�ڰ����&ѱ�_N�K��yԚ�NPb*n/Wk����~�&s�7rFL:⦔�%C�n�T)��J 0��E��5'��jp�������;�:+�:oi'oO���At�j�>�P�1����mv�����Ei��(a2%�2�q���&�%2e�Rxu�������L����ۓ�V �Ra) ��-�^?�d@�dhPw�1(5�"����G�CA��=�G^F��Q�i�;�ϫ �Ɋ��u۶gw�<`��EƁ�\�-L��v��xH�
666���lmmv���#�ҵ��/�?]��GE?�{;:ޮڮԼa���1v�x_���g##�E�3u���3�d���3����S��NBa��;����U�X�3ge��n�p�7O��G��v4�XF�,C>�8�kJ�>��t��t�*����O�h�� �A�w8,��8N���}��g

<������ڮ�����Qp�B��ջJ:�6�D= \��S(hE��<����X���ҍ;���2(耞q�����z"+W6���Y.t�����7����W���#���WG���wM�Ht�[��4;�]��$V?�EM�%.5U�Oc�/�O��G�O���	ݫ��@KS��x�Br��k�M&H}U*56/Hg �I"*�i��-��j�0����& �d�B�f�ٝB��Z�����7��8�B��eI��LX�]�p�#G
��Hr�x|N���a���|�ɺ.���V�L�������8�ܙ,M �2��s�Ȉ��>�F"*��mW
}E0�0�3L�d����]����_���x���e��彲RTD*�-��ۯP���y�b�*zIn�Ar�-,*��A��T��*��軨����;���-�4�p�b	�TG#�;*�4h��q�%w��b�@IC�@ַ���F����� !}�׋��:������i�f�t:z ���p� 2��Y}o��v��{^���CO��*�s�Y<�S��;M�r���r"�˪_��R�����йi50�h&�^ɥ��*�� ����̫0q����1���QYB�����?�ؿ��F�����(I��M�s�"z���TF��L��5��y��-t!����``��<C�d��ͦ��(��}�J�~������ܩ��S���j���#�"������f��/�'+P�^����(Z�`�5��_ԕ��y3�(��8���.xA���f���f�ƨ%!)|S���?��x��~�|�H��r8�'#k'Q��}\����e��O~���ku6P8zq�h0���.��e��`�ȭ�;��R:Tڟ��#3;���Λ��œ���Q��E$���1ಘ�&SKq'�֍@iM�>s��_�cbiI�A0��%	��F=��JI���;@���0 �<���s�<ʫd�iq�h����z��� ���O<�M>}H�Z��ͅ4��R��7X�m�OC*�B����b�c�,=3�]���Lޙɓ6�s������2jh�QZ�*�G2U�zY�J<ژ���b��I��߉��6;��d���|�C�I0�|�ohI�Ȏ\x8��0�oLSB�t�w?/'���������A��@aNU��<�|"��m�`����]؆Q!�g�h�

��6�̩�OS�w������*�F�C��Ƒ:5�(k�u�{�C#Q�g�tA�|��"LMo^����a�7�8A�B���X�v�Eޒ��p9�e���xļ�]�)�yaO�����*&l��Sk�c�K����)�KMU�2<*�����Fv�7�/y?j3#yT���F�IX)XMIs��C�9w�\z�/�_��O��7A��
���Q+ �	�v_���0D�BQ(F�c>_��R���$����֒L�A����-������H2̠��(r�!�0�����*�2@+�ȟ�&�xR��	D���n���X̦�c���H��yh��?>��]��hKfLp�,�I�g(;�q��4��#��a��x~8���N14Y��������0�h@����<w��*۫���UXG;��w�ak�}[�p����)5�v��R�zFFFrK�
�p��HJ�I���<Iڣ�̈́���GGG�cd�DG<�	�\"�Y �@���#E����b�~�:�<�6!+���Xi��477��6��/Ό�L�lT�����(�|C@N��2���M�P�{�$  �Z�ra���2$(ŏ}ļʦf&����G��#�����7���G�v��0��1�]i�	�Ϝ������q��Lv!�o۱b���I�xTxCm�����bxZ�=�	 �h��3������v�d�+�Y���²�����9zh�(Sa�J��RPZϬ�45�˂Kκ�Y�A_ xDlST��B�r�Q0jjj��������5��FX4ĸBWq}�W�gm��[$w����U06�eƨ[�;��7�yR8J��fP؆z�dcK�vc	Oލ�������_^�����f�E,�DE�2��8�ũ8w�ʝ��Cʅ��F+T��|������뗮p�9<pw��y����4MA���vl a�*b��1�gȚ5���!�M@@���	��-ë�������?~b"��ЮҰR�;��o�o���^;0��F����'�m�
Z�ہ�@T�Ә3�+U�v:e;�FO�B�Y�ѽY��/9n�m�.(�yo���:�j,9�Ơ{:�w�.EN�t��?�J�&Z.�� ��\	{%����r�|�p9���&+��d��3�B0{��Ҟ�H��q�f��P���`�����Br}MH�R�οh�3����%C#g���HM����
���g4z��=0���%]ŋ�$��	��&`�˕ٵ3���)�*he
��L[��1��*��i��B�� �#hq��з� �í�^9��)�XO�U�<��9��O5@<�J�6�k�VW\���8ʅ��*��b��dWX�6CJ~���[ב�6/����3dv��ɟ����n{3�4my۞��}����2���ɼ�^!2<�3�V�kpu<+l%)L)M�Q��)u�wX�Y�g�t5���,����	]��|$L6~�Ys��rA+��R2h�E"NU�Poܐ#�~�h�����I�e8���9�L���\��`$�@6���#�b��W��Z����JĀ������DŀQȘ�*Z���ɢ�,s��U��ب%�3�L#�Ή u9���a$^8*jB�@Z`m�Rȓ.���A,�SN���_p�8���@���Mʰ�D.w�/W0)�8��ER�8���>:�6�Q�D�(΍���$�`�\�\]c��?+��L
�/�e{��ƕ���Mo���V6Z��&6a�L�z��X�Y&��_��c��<�؄�O�;pD�ԥ~VӢy�S";B�6���Aƹf�Zǃ�h�<3�ʓ�G�eU;�e�:����c�˲3f��_�5�����#�]GTNҠ����ӊ{�[+�-�����a)����zF�qь�l�Ro�(XBy �띓!��-%��}`�;?1}�43f�9�0;}�Xl�d��!cd5�?�-
M�pCi��F�7?�u�Eo�S�H��p̡/o�Az��*\�$�E��a��m����L�֒�P�2���D�i�š��x��w(=�N�~5��b�ehp A�e��'�v��T��#�~c�W(�BC�3�G����`�2���Vzj3T'6������ۖ��gal��q7Ui8.\��J���$tH`�H�j���
S����T������I����BZ��ُd|]�eŅA�L J�0k���Xf���6CG�S�A� �{�+**�]M�AR|Z!k�Y f�!��Kx�#�#��e�Jd�{6��yKa�> `BC^.%ԛv"�YNg�L�1�my��CIE+a�]Y��䘅ܴ
�z�3�p���-8up�]�E�?������/.���$�F�/�:1ãJl�R�}�U�"�s^,f����_�}pޔy�A~$������ps�Q�
9�!�9G)���b�b���*�g�e5;e*�G�����h���fq�2C�U��Z�H��Ľ]����|�7������~�x�u&���,��  z� R6u�âK����EA#ԫN%^2Nj �Bba<? �C�(�"�����;EC^r},:e�떦��Yv��o���\={�C�-Q/}�-� �m�"����+ACCN�jɡ��Q����`C�-nm1��)Ԋ'cZ#���Rp�c�}ZR�����F���Vj�ML�����!�RW}S���rd�<��C,�%UU�oWm;i�Oj��g�T�I��,�&�%���O����	WR��bȫ@����v�� h��F`�N�s�Z�o�Ѧ˜�t]�0� 1�|:dm`�dE�.)|�J4�o�U��@%�Mg��)K�Aʥ%�^�TJ���م����ƈ��È�P#���r�q��N�/a�*7ʦ@H��:�dƂ�Ӿ8p:�m���<�Nc~���\~,ԑG\������W�B��׹��bV^dƌo[�qHw�l5���m�qg)d�ʓ�چ�v&�u|}V��Xu���w��t6W�~��~�9D���q�H��"0y��]"s�[@�Դ���5Z�K<=+N�:)Sh��`�cf�b�3�(
.�E�TxD�\�'�n�0�o�2l�s���*PfS�ހ}����-�d�K� �}Sd�D4zUG�JN5U�l�]"}�+++ˏ���j�_��d��s�~�c�'R����y�0��u?�B<�_�ur̞j���7;��4��%�`*��n��3l��d��'䒌�q!L'ڙ	-��{?S�ј��_߯�q�he��@��m,U3�:�.̸��q�o(������\�������	RQ���������~�Y��<OH��c��8M�`��Vm��`c�Z�����{��׃xsqޑ�W�}L&��*=��:H�!~��	Ij� ,��H4=K�W�|[�֙�p,6��Sea�`�ܣ$�x8K2��19;��Ty�,۳bP��W���_k����E>��8 Kl�/��,�}9�xhw��K�S����5�W, N�`rT,�"v�ь�O�M�����=��n�z��"�T�MY��AuMw(����,v,�^��.V��q:�~���������M�YY��"͢��G/sm:Md�M%�d4�̿ly�#�ӛ\'�8����0�r.V�W�Qa3(S�U�Ck"�t�����iY~� ���c�:=�>���n�
8��@K�'����ck�k�~j'�d��r��+�OA�>v�K�����qR�k�1��(H����yZ��A�KR�z�o�P�t0��z��U��s��$mv<�AXg)�s��U���� ^�ؾ:h�/�REJs�����
��t�n�����zV��7��U���9i��_�����vm$�	��S�	�˧"�{.; ��`	�̈x����dn��0a4c����w[gb�����b�~�qq�����4F"v��H.f_�0���1 E���V�aמ	�,�����tZ\^Ǆ�2�RbYS��@}�s����~Mz{8�#�ͥC��k������&�9' QRUm
�����}�(L4No���CV�m��J��#���RL <����������Y[��#|Xlmm-M�R�5�i�����n�nov
G��$	�6��ܝɀ��̏�w���Y��#3WHu���l��qUN��Y�?��DH��HF��ҘI2��b�D�6�;��T���j�w۹��6�S	�E��f��,�.H!�AI3�58a�^��#3��#�:�w�	��d�s{� O!�����$Jr;t]q:!^�6Jx
;��b�L�L�%��@��Q#I�)&���H�����j��Nޙ?��6�����8>u]��GyG%=�s�\#�P�uݡn���?�'7�,�ҙ�������%�Xg�@��7��ߑ�0kᧄҁI��?��|~����(GD��\��뷽'�;�C1h��	�?��mSm�{�/�|2��?���^S��p1pþz�6p��/�?L4[[d���g�5�>��_�F�BO�^��poH��!�Xr#p�y���R��D�2���݇�)4���2�f��gӷφėH��	&:��D�ѻ�a�~�dn�ì�|�i�tK��|4��q���	ߵ�K��Иd3D�dvLTVI�XxU��y�|�E�n��W��%����P�J.���&���e$'�Ax L��q��9�!8Sݟ�ʣ �ui�%���xbP`Pg���=u|��cB����ez$��M����u�rs�yDȡ�0��.��'XSn�?c7^&s�D
�y��nAC�Ώ������ɋd$m��_ڪ�w� �W$�" c���M�Zyu��>�+�U���҇���br-�u���dn�F/�͜�6JHo�Tn|�~c��{DZt�[k$Y�v�"�
$�o��z���`��P
�
��!L�]��ǥ��
\
Z�,KU��O�0*�ț -��
�L0#w��{tx�:Dlʓ�����|Ej���:�'Ü9�w��\Ms�ÝP�R�B�M�#C����խ(C2\���hyȟ%_��<~�R]�Q��|�g�0�n���u���<X"=v�v1�;�@��ú�~`>4,�u��>.'H�6E ��#̭읞ka�)��XpQב�)����>?�[�c����?dV�9f,���۷ǸMCX�{�a�}x���В��� l��Pj��Q�٥�,"d;��Ls�'�V�~ڰ�S�gV��LK������Sq����u��vGL���L:�.B;���Gr���9�z0I�CR�J��3`���5��ߌ��D�*,�0=���g^e#{�$uCe[�_E�^I$��4á��Y��8�&��4$����.R�bI�����+rӣ�w3���m�ߪ���}�/�IDG#����m�;�bQ��9��|x�#��F�}��!1&f����%���#j��Gw��V��WEf2%Ś�[$����	-�x�+��U8��|����>eC\�o���-�:❐�6KRxQG܁H���++Q�]��V'���������	6���((R��S��ֆC�6v����6(�0�"��������I֕g��fmk���N�$/�O�e���n*�M� �"8NNZ��D�~�>*hPxq�.�|�DY�m�F6�������N��X��I�8�!��nC �81�U�W@ET�f����ς�^�J}�(ci�L�[u)�X�k^�z�C��+�9p$�<�[9TU��<�Ue�8�1^���X�vV�������Z�t���4�����X�.}%A�aC����5�<�ܽ�"@��#D�'����ޫ̎�WM�n�b��Y�k�A�bZC�F>���1xZiA�/���'$�;��-����=�t��n5���[�HU")��U�'-��^5�"y�r�v���0JŨ�u�/כ$��'��[zP���p���6��_����&ωؾ��g�g�܇�����i�Մ��X�']�Z�α+������OᢺL%��0��0�sE��]UhlM�8ac�%�@�!��0u�Wj����׎O�ڪ̥t��������ͅ�\���<�q]-���i1��燉��4���	�)�6�"��6�V`~ڧ��s���y��SA�*�tq�S	�8у�0�Ⓥ�q�q�=S�[�ё+�T̂��!1t��(0��F�	�����B	#�Y�<����N�ҵ���3�'�Ί:뻲�9�=��1!�^Ab=c��Ī�JR��p��+5�x�P1\�؉x�p���
��q��`���BHh��'e%�A�Uj�mK�|�	sէ������g��z+��%L���گ�� �έ-�VMڷs��G�M4S�/�g�Be�tZ�3�����&����}hQ��t�2�.@*;~�W����F�j�|	3��UaGU&����dm*��F�VsfI�3:�Ր�Unw\��WG�vb�n�7ZiY1�q/�_�����[�Ћ���C��0t
J$+4����{�d`�J�歘3�$�`B5���9�j`�/tR9��wNk��^ �tVzCWj�ܺ��V�2����u����d��?��y˼�Qf^s�ꙋ��ʖ&����I0�����yK��"⬓��G��G�B)���F�J[?M�&
��D��|�4G]Da�����3sG3�/�H&���Sh`�#B�Q׶�ɡ=�I8����;���!B�fde(j��LO��������	4�2��i�S��2&֖[�{P�����=y�*!tc�a<�Q�����B���p~���*ε�ܑ]�O���A�=躻�*JB�Vp�y0��a�H�ag�o*d�uB8�FfU�5�匐��9)�_?<�Rs�&�O�UR���r�ט-4��@w�I8�9ܳ�IZ���B���<t��ͻwU�{"���$�+�o0B�c�Ā'.`#�a��h�f۷�>S���3�d֨�{S���A�v�=��[;N�u�D6�7'�.��~��)q&��	0T��U� h'�*V������m��ٲ����2���4��!B]*���Z6�gD�>�bGL8v��ް�tP��G���)��[���N�+p�U#��j$G��{J=��.�[5�i!0ѓ)ˉ}AQoK����o�l�ۣ&�c�o#���w�����f��� �n3�]^�n1
S4R̕bz�P�w/f
�P{��i�vfZl���F�)R^dnb���̩�zO�Zk2�
W� =�4<�	y�d�}�O��Tm�W������𦶼���A��m5JH[��/5��'����H�+L�3���9=a���U�-�^G��C��γ�5��$�6�pl��Eda��A�N�F��j��ӝ<�𭺑E$DAlwyoL�]Ӹ�"8'q0Id�+��\�����Q�CQEt�\i/m�p+�e�,�Q��*k���_Ȓ <����|}Iu����R{or��!����J��g�c�h�>S�e|�O��Q(<��R̽D��zL��H�nۅڱ�2�t�LX;�%?Q���'�R�m{ˆ\<I|q����wl���v�о4y�'f��v9� i_ս��ƀ��Nٜ2����p,�SkL��x~�5T*/�hq��ټ �T*kT67����#��������V���[��l��bN�)���#FQ�8�O@�ֲ0�`�+��Y,��X� //V��/$����{6�~h��j�}4�l�A�t�7�T��`Ug��ZXҤ��H)�h%�5m�tI��v��ƞ�0[@��n��ބ�$�^��,,�ǲ`S��~�t�z��!y?�X��⽩���GU.�R��&��h������4���=��=���.���.S�[dr���@˗��m�\ʱ�[t`�e=fPl_�����d���G���S���#�~P�D���ݻ��%?�L6�����9���q���׵�e��(��j�`�|�:XUNLf����.�/����|CĮ��ვ/��;�L����N ��%�V��f5G�Q�x�;~sV��
�i�[$��r1?���ߗ�����0�K@ް`D�ϔ������ ��WR�zb��;���*�c��Ъ(p���t��܈D�Y�����)G��<�,�=�B�j�ӘыBk����(�>UR�O&�8v�%z�F�N]up�)��]�΢ń*7�J���\���J��ԴI����'n�s�)�_�D�
s�3��C�#��;UU�rI*��庘���q��4� ���^����U|��W�-�co�@��)c��-�G�¡bgE�<��D�ʫ:!\7`$�$�S���ȋ`101asA���}�(�A��n
�5�6��J�S�Od��ak�su��d�]	1�]�%~�b�+F�zJZkߧQ���z��&�lM�>+>v'�������݀K������S�[��5>5s���o1�ʦ��}w��aѳ��o*)��G�!�]e�"�<�]U�� %[NJ��/�\*�?����|��ן���IC�&�&���+;�����C��w��@-����-�.���:")�R��������9��Gtw #����9jH�c'�� ��Ic5�Ve���/]z�xP�9s��P,�%����F��/>H��P�3_�܁�����s���B��l��ˇE��{�ŃgdW��F�S��=g������S���y�X�z�И.���d�N([���SYt�#�˺�ӥ��æ�w%H�j��-(�[�-b���oZG�oE�iYf�3��18�� �MYN_.�P��%��{g���=����қ�21���O>�J��)�׆��;�z̲�Mp)��f}u�ݸn����ic��A����y�e��}� Z  ��F�����A��S�t�l�}���ч���iD cm~�5_?{�/���R-3,hQP�ĥ�`S]�E�GjGk����R�7ӎ&˷��O�P��}& |3 ����]T�5t�^<V�x�J�sh��}�ߕ�@�I_\��	J>'��I8�ͬ���i�T�:t��9��GO��ad���������Uָ�x�%�P�gd�We��-���&�����E�H)f[U��<�8�T�`�Y�V�Y����C*��eΈ^S�� �SuLȓ�������c��2=�O�G�����Ds������؉c�5�����Qq����גa}�-�"��1��V`UXQ{,�M�WO�����:'e��#�.Z,8��C�~�5��<-�E}�S�Jdy�J#��<��d-��M���23#""�F�(U�dU�5�t�y�$(l�5k��>�[�1W2GQ��	���[D���}�7�R�0b]�՜"�D�;�rH�a���A�$�ᮓ���&MV@� [����{�I�eƺ��A�i��W8���<:�������חB
���r�	�*2˖��L���.X��	��8������Ñ�F�I�ҥ��q��G��a��A�Ѫ�,Gu�}��	�,-F��'
�ň`�6�/WTD=[o'[�x��U� &����vN���A�D��AՇ��f�J�f$�y��?���yj�I���Q�C�p���̒Z��4d�B�I�	�r�zo���i��u��̺�R������R1���>�9��N��Q̰�h/`��\��-c��E�,_�� �YRp	��8���84T�_�Z����`�w��&\���B	��ޯ����<a5�/^����Nka�i���[�aI��b�@}%\đH�7 �݇7L(	Ne-����e�o� �XvUu/�~�_��'}
xc',����y��Xb�4�b���U�Q�}���B�4�Ѐ��.�?s6Wu�scg�97e�O2�;�g!�!9�5�ɿD�&��H���Ҡ�N�����R�m��8b��*Ӣ#�,����[	�cA���J��O��oއd��f��]M˥ sۑ.�-��Pq7��e
Y����H���w���3������?ۅ`�`f�5��o��Ҙ ��#�J�}�ďS�$�I�(�F�e'Y.m�̲�r�t2#v7J�eivC!Cz�0RHd���Ch�
%C�Ǉ ���K�O*ҕ�79!��A�聢9w���))i�0 ��^�$�gxQ{��h����zoC�
fx�9*r���t	&�`��܏]�W_��a�m���4��*k=���Q1�aC+	�Pw�{�ӎq�֍��Q*z{���D3�������W�-��Jatjs	�k����Fs�Md���߁a$>"D��&�@L'��;����"���	�����	�%��C)vsC|X����S�O	25��>A������D���"%ty@:��*�k���|��J��?�yw�;ײ��O�jǵl�@����w���Y�c�y���,fV�����}
:w���<B6ꤠ�����3�T�l�ЊB�N:*P��;5����C���������D'B^�.�ȕ����8L�Y��V���S�����$2����N�溳��q&u痭�}��MƢ�ifS>J�����ٞQ�w�w���t�^{cߥs��tk����$���
���@�ǈ����x�b�Y����1厖�>q�Q�I�AG��RQv�o�p�J���$��F'v��W#5�\#s����	e�"�f*�r	�K�tsӐ�>�����V��H�HT����^T��_Rps���f��J-��IB�qtAkiWtnD�_��UG�N��4��F�z��H---��	��秧Jy�44#�E%�q�ဘ���)8}:�|� ��(������\�ϙ��[�q�SdJB�P��V�-�p���G_<;,����F�$�X�i����_̊�����j��L�eu1��"Z�J��zX��¼z��#�xhMl��8Z٣d�Rhe����d҃�!�� (���ؖ�����Z1|�kh�,��-ZzF{̸���h�$h�-��/ۮ����N�G�-���r�
�
hJ5����� �I�e+�6��7)��2�Dy�B֞���!��'x�:�+-�$��fG���O	(����y��A;^���ޘ)��K;|�����33�����V-2��<����_O�-J5P2��4.�ł<n[l<8b�bK�Y����$/�E7?�|��%�*��Iђ�P3w��1�l�X\���IqK��w$.u����B��3[b�!���{�-��)Nv�fs�9��|&�%�8�C&ŋ�?���W{���3�\��:gx;��%۩��g�����{��p5���I����t �Ƌ���������vQ2�I�_��Ì�/�����Cj�o���*�j����6��Q�Z��(4��)�4�����6���:��>�]��؏s2j<��FEH��&�b�i-f#�B�С����PU]�^�x!|�ܵE6F�y{1yq:�BXBg����1S�#߆�ף�����K4��%>�DS�h�uЙ��ig r�W
G �<����
���_��!\�j�ۗ%�hrɧx� kk�� �jjw{�"�7%ߦ��C3�Eh��t�=���c�O��s�-p��u�m����Y����,����Ø"��6F&S�Wk���JbR]��|��Dm�!�N���ַ��BJ�����L@;�Y�fJ���ӆ����|]��-���k\�f(�]&�*Zy�8�]���*�uȫ����"Ő�K`}쵯�AAYJ�8�NLSz�'��B��U������ގ�U�-$o�rFWY�O5-?�F�c���n���?��ֶ2��%|���w�`�z�<�^�)V�.2�L�/�ѻ�w=�����pZ@{�<�<�깉���R��x�2���i�Z;�I;Y�m9_2��F;���3��,��=;��_Nϐ�5���>��]As9�ٽ\N��+{6!C�_��3٫m4$��;�>3�zw���C�Em.mծ��QB��Y�-v��`*<l�����n|�>����Z�n�����d`y���|�{�t��O��0��W�f����gc���\H��Ha���F,n4~��]/_?AQ�o!�'ʠT������7}t���~n���mkd��	���cʠ�Y����C1stS�rG\�k�^�J���.�5?�@DE�dp(��muF%����N�
�$�GWr��B�Be;V��D��Z�G'�7���ʑ�;ל���b�녻ùW:$��EJ�P&J5���ZYBK�Of����|�����$K���!I�t>�|L�Am���3���5i�)� e�sy�|a�a_�W����ۗ��V�ԝ#�c���� �O�:�r<�n���A�n-���8ؽ���{��K.NOy���V�kǸ��r�95��V5@W���Z�\�w�gE��
2�A�#�>���o'�#&ʸ@��k�T���TUe4��ʚ��3����(��@'3�FT��MG�"��"�^�!o��I���0
.�`�	j��"����Vk���,1�4T\G���

>�7L��[*�
�U��ڱY���Q�>�$?g`^N�f���a-(�5��3[3���s��u>�ܖ�^�u>g�[�|�ha;mϻ:^^@����j���$�Z�z�BB��sħB{�H�D��/�?��ä�{4�K�k�^*��j�c�U�;��JN
/��@�|I!�G��k�����^Pg��s�L�?nO�抂M�8^�����9��eW{[4�bS�nf��e���C�ҵ������~I��7e�����\a���x,���,o>c�뿑\'��N�a,�#Ek�|mN�R�'j)��M�Un�� ���:���m���ۍ%��q=�%�����g��L����� ۙ��o������`R�5TL����O��f+��`��������tA�T�Y��y�����X=��mm�]l���>�/{�_1��i����	��Pk�z	y���kϓ����瞓V44�y|�a�5ק�)�ĢLމ~��僬��ӓ���ˡ�� r`��
Д��b6��y�q5�������"721���F�&������n��C��޺Ӕ��Hk�-%r���/���/o�9B����16K�[v�~�}�
SȥY!�g��Yd�Z�r3�5ⶪ.O)��m��dt��>���@"�Ef�);s��쌛�m]:��qRZJ�8L����I7*%yc���m�0W6�u��9�&�⺙�����31�^��%`˘!�J�Pϵ����4mx���+%}�����υ_iR����,�|����C��L+�c��_fʃ�|���5�w1Q�X�ö��P7^�}�<���G���@�T����c�묻/��>��O�������7��g=�� �>��7��6��931�v}��>#��ar�c!k��nW�c*��yG�<^�637Í��}�'>U5Vb�Xc O�Ҿ��`:�$����[u�s�Y���(��u����߱PP}�%�B�,X���~"�n�cZ�yb��7Uޕ��q~.ϿŧzmG��Ƃ\�]��z��T5Ā��mBo���d�ua��t�h��ʹ�(܀|�?wa��&,6a���H�m�u�ߴ_�S�֊S��{X\=�\3]�
8�<=������^�,7pɋ���� V(M�E� :�:Cz�x��+=J@��@� �maF��̥������5g4p�D1'��f[r����x����P���v���5a�~��<]&�絠O��_=���z�+���������Q�!A[ڥأ��;6���D@{*d��Ĥ`�6-\��������_�t�kn�����
���.[e��Y�Pf!]e;q�Y����;dtV��Y�9{�r�	Q2��e�p����}�������������EXT������2T����aZ9Jf 1���S��R��+��n�Nk�es��:�A��A�־��ĂP��tL������|��N�(�̸r��,�`nf��m��q�%����} �M6ϫ�n��[�{��eH���u\]�����]�@�S��^-��ʣٍ-N�wv}�R��Ƈ�Fꈟ�t2��+G�~5�����)��lWcsm�i-������,>'��t~����2���ta�i^�a-��XO�)�c�]{=�c&$�*ݢ�O#lĞ_82���E�KV�e
��u��}	T�y݅�2�u}�q���{�9�r�Pa���{��x/�c�wH��ַe<��̭*���%�-�w���/?�,W �O�9����߳��K?\� Y�[KM[5�Ty���C��¨�Vs���l�~��E�<�}���~{����~S	>6���G�VUŶB��N�&�lh2;��دHi�����!�-)�f�����n���Q0w�(�z����FZ;�����QD��Я�z[��H9����a��'��e���K��	L�G��{�g��)B	�;�0_iF4�(�ab�'�B�9W]~Js�����x��]B����t���1tH%Z��}��eq/�;��Uc
jW���Dd���R��<N�c.�,���s��P8��-v;/��1�
l뿨� �Ok���ܬ?���ޕ�>�	q���G_�4͎|�ѷ��7�*5x>��?V'��/�8��5��<st�.��*]��Rr�~��������<�Z������L^h�.i�<��F�@ m8mr0�kn���̝���B93��Ks���_�~T-s��sj)I�M��s�3�y��9�Q��V�\��=G������D�Gt2�Պd.ǭ\GT��M�6K�fT멭x�mTx-��/@�2�ظ��0R^�T�zr�Ѵ+/6��*TЇ���R��"�X�݋�ẖ&���G��Jj�)��X���;b� ^�ؾ1c�=F�#��W�D��tH���w0��4����l�Q�#�^���̾.�_��p�z0�O<ϧ"�����B�׋�3猭�N�V�{�ac�uF�z׳���X9�Uf���.S{^��aDR�;.��O��i%ϴɋ(�	o���{�~�-���룳%A��%��&�=���վ��N{���~�:d����yd�)�*��mĥe��k��rz�~S?߉���V�?�P[z푖�ˁ �i�2�o���PY~L�1O�;�8Ja�����4Lw����/�t���[cɐ��5>�'�b�z��!�#k��Ƒ�`��#��
���¶	�[D���}�� �S�O;�f�E�k�I�2i��1kJ��W��0'%r�	�%���Z4p5jH���?ЇLe4����ic����.\s����ՂZ)I'�j�1�Ws!�fbKTJΥ{
�7r��{���X�o�v9�~�]p��.
-c�׎3M���Uٳ��eg�ϸD+���'�ٚ�,)���ɧG��+3zxHD�j��IOj�\�tR�<����L]Kc#�
��I����o�.�E���b�c.jm!V�� �K�[x�F%g� t��V�Ja�����?&���ȯY�Ώc���O�M!��B���(
.���L
ț������n-+Η��C�f�O)5֘��Ԋ$�����B���X�qe&!��X)t�����m=Kh�7�'~S"�,��Q�9����^5q���Z���!w����S�4,̅,^h�uE�8�~<%1E��҂��R����R\2���ZEL9������7�K��r�w�6F���5���8�C�6c5 F���9� F�,����ZW�}`���VUU�;�	�):�ހJ����9��i���M?p P�y$�
�O�^y�����y��#��"�x@E��`�D�U��ȯ,�L��]i���h8�p���g�DWYR\�-l��p����|��oh���&�Xs�QL-�4z�W�[hM�J�0◢�{��g:O������e]d%&�\W{6.�_�!L��;��g�� Yc�J叉�4�;�4؋d-2��i�͐�ng�9��XO�H�W���mZ�Ŝ��$�0/2z1Ñ7�T<�k��M��t��k��dR��ٱ���U�е�L^s����Lf���F����U
G����rɜ��^�A�2��{4�ps]����~����l�ᷱ����߹�������[zA�u<�)B���֮���'z圛�97�Z$���/:W���������0e�&�DN|�����_l(vt�+(�U!���^������{��Zz���¯��o�c�F��q���;i*�O�"� �z{�Q~�}?Y�������	��]U�|ņ�jpȫ�����º���&��Fތ{�@�,C��۱��͔�G������Z�c�	$����D�C}}��U�ph�ִ�P��q-T|T�^ԧ|���B�w9e�;�\��U�H:;�1�닧2-���է���q�K�2�nnO�����PoS�3�P��Y�D�vp��-n������v���Z��DSQ�8e �`�G�^
�}�nt�>o�+��Y� )Sz��;ar�#	�ݸUnHs�4�uڧ��ᏟIs��N�/	C��r&:"]���)��Lй!*wQ���*���\|B�O�<vd|���r�d9ܤ�1��"Wz���eXh�����˓YY*��Y%c�M�=��:?�ȏks�{LI�%f���W��G/D|�q��+B��C&�ך� Nj�_Sb�+�
.HS+&�T.��Tb�(��
�5ns�ν��%�>u��ܸQ�8�8�r½���^߭6N�k|N�މ�m��B��Fz\Q��צ(a�%�GPV{A1��2O���s���
p�i{�)�9	{��8.R�x����.���;�m�nV� ߑ�
`��1m��]����YZ!�@L��ݬX"�5b��V!�H��!����"��`]s�#	7�<8ٴ���?<Agۓ�w��lkA���Ag���i�Ǫ��D���+d/խ�����*L��%@�v�p��qA�_�t���5m��PK   ���X$�8�l  �  /   images/aa130aff-16e6-4627-9689-819d55b5861f.png�YUL
��Xq-EY܊����K���a�RtY�_����;��kq}����M2s�9�L2�3�/Z��X�XHHH��Jr�h��[0��Ÿxl���d������?�m����p���d��e�j�����e������ي���&�D�	�F_YN����3�z����k����Ԏ����(�Gǳ��R��7���c�JMNf������a�\w��{�I���kD�b�K@�)u+h��,?I9=̚;�����[�(6-�r�d��CGG�%��+��1A������G �����B���	�A�eF,M��Lo���k�=�8%_<�3��5���K4�AlaA��~��V����6�~nU���٤�:Ƌ]��d*
����W��CMy(%.KL�)�U~3"`��&���Y�t t�I� �Be���qkP��r�<f|0$L(��-+_�a�� m���$�J&�a���%���}$?�}}����4��ۏ��˜
|<gX��m�/���&�f27��+F�lȏf�{L�4d
�"��)"eN��_���`��N� �W��ܥ��d
ڵ��Ϳ:��-�^���X*�^�☈"G��oւ��^���i2���n	�ii��}I� ��M�L_�n
k|��g�^�D���Fg�Y�U��'�Ԥ��������$k_{���A��G�1�F\���uGLvaf��<V��W��f^���2=Wt���\C<�m&�	@�Z�O���g4��͆R����թ�#�7�Ȇ�A&��f�vf5
�"����0��hż_�z�@o*���I�3Mu�l#�c
���H�Z�I�C3n���6���ﴪ�	�,�@_�7���E_��~��ܫ�[&�N4�X��������'I��^��D��;�d C�uI'��;�����L��ږ��!�@7�<�^�����	�ʉ��!Zv�pt6�L(�QbG���Y��XHZ�e�<Z�L�$��K�V�jN]��{��i[E3<ӿ����R¼�`�ӡs@^��pv�Z�#�A��4d!~�D��޳%�{����i)�*7�CՐ��\,��{�_{A���>�Mu]hm�w�bD!�$_`�12Ő�Y�D	�,��&���W;��uo��oX���N��������c����`j������{���c�sH8�0'ޠ<C�ȲL�Q�ۗy�ߡ`��#��Q� ��y��IX��L�J�{�X3�̓0�1�|'��f�9�CC�U{�'T�K�c0�W�&O�BMJ�7&�꠰l�j��������X.7��k���leY#zu9`�4;��w�}U�@�l�`V�[�Zl|D`�eJm�c嶚��lnQ|l��;�l-��|�8�Z�-b�P˪W3��OIƭq�:��KS��d�iؤ�)��)hDסQ����UU��e�K��iKR��@�^9���� ���7G��*�p6�����Ir����1�q3��	
�Fl�I�=m�h	� }9!��m�W�:�1�jC�����w�(��b�������l7��2�~xJ�֛}���F\��w.5��ߔ�h)UV|il��;��cL�{K��ty��{ �``���C��p�w�kz�����I��g�'y�h=;�@�D�{:j^.�m⅊��|Ǚ9����;R�ȍ�� 3����xw\���CTl�y�,u�v�e����Y�(Tc4@X�l?��%:��v�M�(��� 8�TZ6�[��_��Rz�#�E)��i�{�5��.�X�uj}\m�w��~&�e/���H�8���Q�/���H�R��5���_�5�q��i�V��;���~�++�9Q����9=�CK�;G�T�N��㥲b�=;�p��>�3���W��.1���E�����|��Kv4/�t��XTJ��6�u{��%Ǻҟ.���G@���:� ��y%��
��E�N7(�� 2�-���]�H���Z�  O3�*韭�<m\�����t�pz�#�����Ց��Um���C�nĮ�$�e����uesM�����?����pc"a�4u�hi� L���(|�ϯI�L� f'�E"��*٩��ծ� 9�-]�]�������S�;iSKn`Uȏ�=����R��8�b�96K�A�E8�կD�h�⢛ns�/4��b�#5���6�R^&h`�j�y�9w�T��ێ�Gy�x˞�iz
z箹�c�*�_�9��Rg��U]���,.V�m
g�H ��rK[}����цQ�I��X�H�����rZ�y~ 
�6M��
򗢧���A7��!ܡ1�@��I�ĩ`!�j}���%h�	Hm=M��ğ2�2���I	��F��[�!�Myv�LE)v��� 3���>�xj�+�Ҹ��_��a^�h�$�ՖL����q�Rf�.��� ~D��O(h7G#�<qF�[)�������k�mFG7fL�o��k�1ջK����r�W��o���2Q	-��k�z�Phiѕ��"0����u��{���blRxk\�SK�.wFM=gx�)���;��(DCR���=���}���ST�P؜f���M��9M��X��Jlָ�.�1Bf�b�^�����g���H��(�_��_���	�F�(�P��}�y�&(�$՜D�Կ!u�y����e��a��,2�R;���ٯ��=����"3[	���6�rm�E?\L#vO0Q�3g��ˁ��m93X��GS�=]��F7/�=6��z�|�y��0�7�#�����7�}m���4t��`���H�袟���P�N�ɖ��{[���4xʨaO�K3\�qd`��R��sL$����;QE�I��G)o�LQ�uz+v׺,��L��X����%�\��p34p��Ѩ5 �j��Z��g�<6�^ܘ��岓d$^I�@//�!R}�V2qPN��H��b5~�q�@ ��>Jɒ��3��?9��yb�Yř��s���1]%���Pf���&O��O�X�����S���cܹlb��Ya��@E>��7X>�J,#�В��s�*.i�JeyL�P��N���	�@׾q��/"�M�))��u�:�����T؃ZV&���b��(��h5�]�+��9��0�Y`/��|�~�<�����d+�_?{����@�U��bꎘ�״$�P�`oP��R`]���;1�9<P���Ιd��`��rCF"���\ջ�(d>�M%DiJ+(63�Cb|"&��x�xL2%ѼZ����CV(�(�aW`��m��R�E�o�j�SX�r$�h�cz@�S��.������/���kW��z��[���z�K[�tK�f(��z�ôڛ�I�����r��,�*$��;$�|�q���zw���ǜMh =J�"2�Ƥ7���"Q6�˪]p̻�Aզ�s��:�C����w�5�hxa8B�L��n{�?���(�͸nu�$��Lt�z-=
>�EO��M� =�=�pΆ�0٠��Q��e�Q����_����h9>�Q�?O$W�d��/?-��uh�4���)(v�Uh��CJ���/Y+���<�!�Uw�~]PP�����Qǟ:�Ǟu��o0��|j�sv�%�U�d16͉-���Ze��Z�PR�_Y���7�������}���؆X����Q�������)6�	��N*.)>�.�G{��3�L^�u��p)��ÔA�Q��yM����Vp,}(Ll�xh�����---l�PT�ruru�ޥ2c:��n.1�N�\�4�M��3�ť�N,��f�e�����5i�@�Aɭ�-YQ�S���fƎz�
�*w�ÌO�ƪ�����'�J�/���#�%��.���U/��G�+;�ET|VP8�FBM����k�WY"���>ފ�]Rl2�T'�w���QK~���O���҃��b�15fBv���tA��g�q�<QӳRolև̅����A�D�.`7����B���*��R��$�ka]|o[d��J�=Q7�FbnO��I7#b�F���3�|�T�#1��D:��/MV�u��Be������u8T��'�&*�c��/C��̊�|b���,5|%���l�W�d�_���V�{������)���y��4C�dZ s���NX9�[T�W�⍪��ѵ� �"*SPÅ+W!��q#���[Z?��Vl���{�w���	�h�i6�XJ�/��I�\#�)짎��~��x����@�'^�u�! "F}���P�����@f�kM���������`mO��3���((��MƠ5g������본��N��_�b�mjВ��W�O�٩�7W�}I�.N���وa�lF���ʔG���N�$so��]�S�ee���=~뤶��@��N�z�5��:�s���ĕ����R���5֣o���laӗ0���>��^q�������3��2��R�7�$�;;M,ˈ����B�������`��W�p\4�\�qH��� `����1�T)!ؒ�Ak�J��b]��%{���DW$����~ս��F`(��ÑuCg��F�(�+g}}��'��- A��x���6����n���#<�]��a�������{�c��J�,�5�p��qp#��R�ZX�S�/.t�Zr�]A��a�N�(6���_km�mR�c$�<Qq��)~�+���f�Z*pk��Z�f�͞Ff�/eꝻ!Z�@�`ḋ,����?)�*��(�<E"�3/���"���"��o�{�RX�N��/�a��ZU���xm��iX21�:1}�,aS缈M�rwg�xM�u��k�Ѯ��e�k��V���S�Y2�֯�Tw������o���];��nf�/��ŧ�A��\��W�o�@��sފ�H�#��3��m��{"�E�Ӛ�G_�U�]��K�i�,�E���6��tl��$N�J�%9��{�P#6��䓏�#��.�^YSx��WBI���7m��O99.UϹ~!�t������	�[z~� SX]�"{��#���7��4w�M��z���$�o�,lM��u�D�Q���=429~� �����AŚ��Zo�Fc|��a>Bz��
?�.j}�"�F�4�'OdZ-�QB����j�IF���{$��dֵ~�l�EV&y�˩ XXy��DJ��c��_(}��s�T��Ҕ��[��D����Mfod��%������Y��cZ\���$�1�\�Tgp�ڊ��-��I��*p8�C��k��Sm6\�������<� qN�&,&L��0���=��M*�+Nol�X�V�ډ���b΂��z�o�����ӭ�������YĶ��U$��H��)�5�:eW���Z���<��c&j�0�b�m�վ�s���X�O�0!R+"����U%���a��b)�[����z5g��x�$����Ke�����d�@HN����c�܂ח��):__8�$���8�+�Y����JG�짽�4�E�^y��5p\���h��VU٥���h�븏����|��^����ЉO�I5'�V�t=`�},R*G���8Z�]��Bg�X8�F!�E�����t���2;ę����+ݘ�V��L�Cc}����)[�-�� .KfwG���<8^h@`!;��6ͮΒ��z�Z�%݆W�Z>;�[��#���0�%�o~���<;z5D�)a-��X߼}��U����[��̸��W>[��
���D&yY��~�}���cx�3��Ey�1�VC����wv�Ӝ�)1���Ⱦ��L=���V}8�LRo��N� <���5���w��x�4����O�߆��Hc���]H�Z	Qi�{�������ɳG�լٲJ�����̸�V4�$E�2�z�5�|�R�$5R�a�qL�qe��"V������X��	�y_6�IG�41��n����@l"�oz�i�v�ɤ��KlP�*$La��B��g4��i��/��<�:�\]/����d�!`7��k��J�AVf�����Pmܠm�g\|����"݇�P�B�?� �jdԇ�-�#u=
n��m9/.��\����\�]��g5<�����y4�#F��C!;I�@&0S#��T}���wd�@C��{�K�H1��7��,���M/�K>���-N<�6��"�wqN�5���s)��G�q*%���9L�Q��0�wk��w���x>0.A$���-�?�˙6/�PDH���>��2�P����Eiap�13.�U�Yz�C�)|�s�VkV����#(V�ʹK7�������ߗ3S��n��?�p���gҏ8��Bقo�'j���BbZ�%��M;#w�"�⮣c5~���/��IseIu�/�}�m14ƷS��b�#�<��k"Vj�͇�[���V�o묆I��?DoA	�Sv��&��������d�~����6��v��h��=�X�?mΜ��k{�����6�c���W�L}c�w�.�S�~�Y�s�_ٴF�u��;��8���g�����QT�0�ap2�;Z�1''����>���˵X�D�%!�$�ʽc��V�/&^+lB��IJ�(��y;����+<���V�ܮ����z���Evu:��2����=���!�K�[�xWK
�il�����qn��>I���-��UI�rub�j�=Qut9�{̝�#� Y���r��q}�V����� q�n��6f������O������e�� �b����`���g��8t��A�ש�x)n%�W�7'��C]$�3�������M�s���-|��f��9��A4K�l��@F���D�����,��ߜA��[/"*����%�="5=�He;�^	1#F�,"�e���Zo�^?TV����_��z�^ЦE>@�
>�$�RtF��1~vu>'��s��K��Wk�pϚq���A?\7�~ϟ�_�G!
����&h4�[���

d�.����g+�񿩧z�N �C+�ޛoxt��mS�j�����;�'���kpڜ�L�]��)V3�� ���R"�@(����l��t�O�;���;�
Yͣ>*'�a^9&۫]�g�7p�v��W�&�C����C�ޮ�����lloP�H�l���(�����X����}�`���cZ��S���h݋�e�9Am3�P�<(�L��ho�|�h.Ϲ�о'C���F�"�ʉ苃��7�Jpk�xsJ�3I�U�X��V�D���6 �OfQ)R�R������r�l�i��Q�u�)��-�a�5���D{j�b���5{f����컈@����㠸.;����}l���p~�;(�:�6���,�y��{?%�9민
�8=*��I�)is��c{�{�#diۥ��,��lhq���W�!��a s��[q������%�U�?J(e(�T�sZ�%�����>��RnӺ��j�ܿPs�>��l��n�wEl1�u��O�!D�	B��Z���bC�~�3Px0{�#�PR�_�L^��,����A�ǁG�	�?S�א+}�PK   ���X'�Sz�  m  /   images/b4b7fff7-3733-43f9-86f3-7eaab1c92eea.png�WWP�E �$�.��(U��TAz/�J�.AzI(FRT:"A@� ����P�j�b@�����>���93;g��즚�2�x@  �Y_O�좺_���"�\� ^`��m p����ma~r�ޱ	5�E�{ P(����o��K��L@���-u �対�-��|r0�����|{22SԈm�����J0��d�]��r�2�~�:>������OT��9tW���,&Z��IB)����Me�iQﭹ/��G�����vѩ�6J	{NԜ��O��:(s$|�T��a�k�W�jjn�cX��e�!|�1��/><=�Q�����uu	Z��y˜��{����Z�xc��8ЮP!�Pݏ����]��J�x�nUz��tY�KD[N/�!�n!h�t�-�)�ZT����HXQھb���3f����cn��r��:����?L����m�?����#"�_B>������+ń�N�O�	'�a�!S̡�ɳ.?�K�+糮_�1zU.D��R��s��LM>������IZ�Uy��N�ʻZ�=^1����&��/�j�{~�B�6�$.��h�	b���K�
�Nv�5<�5U:�ش��ґ��]|dӏ`U�]g9N+`��&\g#�&0Ii�~Wi��qF��G��Z�ɻ�<��=F#P��{�q �?�(/M�fś��&����ؖ@��9�C�L�r�KV�%���gV3)"�r���9���A�1��K����&�̑~G�ZS��`����z�@������2\c�)��u���fY�U���J��������t����N§��r��n�DT�ם��I�4ca{�4�R�/g^�Z΀����*�]����6��H����4�����ђchw�n��In�9�6s�kž���s�_�q*�8lJl�$�B��J�^!���g��YGTW��{�Y�Kv@�~C��N��p������:F�I$�y/���=��}e���!7	a�y_�,D!����\~��G���1K���۽��P�1�^���K��]/��gi:)/DT��ձ�W��4�e�����׻�TP���N�Ĵ�{�|�~+� ȿ��TfT��_v�]z6\4�^�(�/�?+r�^�-�R\+�d�߮��`vͫ��I����R�2���#�:���\���/����2~�ޞ�6�OT��A+��U4 �{��V�n�L�9]	&u�Ê�ʁq�c�IW7F���&�ڿ����:�}؆��٣��C�ܚԟ[k�&��>4/irƛ#r;���?��!�:�Q�n��j��p<�@B�0�?��`tty�j��~�✫~����]�͡����}�`洴z�hw�S@'2f  ��!=�7��r�\�pW�쨏����C�����xI�����TIΨ���Q
B��������������D٘!��|�^���t/v��_��M�����-9
�ںmE�m�K�
��{�(��yw��2'�y�4)K�	�WN�4{~G�"��p�^T��W��z\O�g�Җ��N��?��g�g�a6j������o{��xq�VD���r<Q�R�.Fw�����X5�͑�wQ�d�@�ݕ�0(�!`�5�6�8�.HלI96�<��X*����AoV��W_������ɼ|����.$��ڎi���J��Σ��j?��1��Ս��tƛ�|�;N1b��3c	e�~ͭ�W3ɾ9�2	4�';+�~1?מ�\np�E���@�9���4��V	b[>tҗ�Ψ�\n�O�G���B�$�ܯ��l����bH���r�(kDJ��o��������50qu%�Q&�l��q
ah��B$@��T�>3�=�KR�a|D,�'�RD�7[w��p�e�	m�`#6�-�z��/�R��I�A�S�ݥ6������H�G������׸�<Ի�}͒A��)��?iS'۹�dq�@0�p���s�uD�EJ�~=��[����\���Ű�˺U�Q�>�N=�)ߡ��h����Q�C�t�V�g4���5".TkN�l[���?`�z �"�����9�� ;41�r�0Zv��͝�9��E����hth��kK��iea�a'v�/IT����"�R�aQ�2��Z7�M�(�@�8qf<	҉x;W�+�\l����?��߫�å��^-MW��<������:�[��(�Q���h��6@�2zP]A<,��3���F��[��~��6͂�J>
өQ�Лw��z����	8��/���M�W�n�=�ѩ鮎(�O��N���'�bSK���%��C�L��M*sޞ�嚖?Js6�.Hz#�o`�]�k��Ӑ�J�}�gA������N��[��j�
���&�u�Z���,4K�:&��V����W�����w����'dӧT(��ϏvpI�1"���ԥ�[�N�C����l^!����d��[N�\�������y7�s�������!/�B�'S筱d��(
�f�Lc�� �ϕVG�֜�y����Y�W=X���C=O�x�?�}�Ͼ�T8Ab���'�r�}����+n����o�8�n���Q�8M�ubC��S-Wׇ��Y�Y�^h��K�[���y'�>0B

�U�d��� �.Eo���v�[W���
��mYe��>=Gc�ְ�36ꍽ�J=�U1eR�ѲoR5�q�DL���>.o�ps���t��&�V$�P���s��H�3s����t���kJw�Ɠ �K��YK'}4�����N�; n������`��~�Py��S>�_}�ff���{-��h�YwaPg���UAt����#�c@A�τA�5G`��{� �'an�')�,�8��&���2�>*BaW�c�C�t�5�0m�niz���M�c��I�0+�Ԭ֢7��q��H��d;�s�~��q� ������83�{�h/�#��nC��H�߳���v��M.�����l�ýM����,{�	�!b:@��LN`�gIZ�I���]�MK��͚o�/ܨu?�Sj��Wbo�	���ԠJ�1/f�S|����ۆ����VL�
��d'�ߩ�y��
��:n�P&)����fb ����T��>�W�Ŋp�/��>��R긥��O�9���W�J�W;�Nff��^8%�Ƿ��R%Ґ��&�YBi��3����a�����r{t?�)��⺜�D>��avN9��/:G�
]���i�alMzy唣���>2=v��"�DD����MG8�IYfڑ@:��?X�:��[t�<�MT��h�v#�lk�.��k��j�i79N�n-N�Չ@�ۇ��%
���!ˇ��&�M�i`,���/���;q�t�쩉�%��v���^���`5��o�½���gnΓ���W��������5������+ŗ#S�k�#�g,=(�.o��?~�8�~PdbM��z�S�Q���i�v�o�ք#���Y|�n���xSS)P��Kq�1��J0D����[Z��u`��Gmo�$}�:����8	y�;���7{�?Lg�w[��w������__��;�1A���M|��gJ$[ܣ��w��{��M��&�-VL�FB@�L������5��_/D��{9�|e��\�s�i|mx�S��9i��X�z���R��%�sہ� �1�l�]��5�^� ����ɲ�5Y9�9�M�G�V�׹�{����Yc���7i#���T�S���Ų?�D��^�ˌ{>~�!��82T�;����ਊecС��D�S���W��X��L�/PK   ���X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   ���X���]  [  /   images/cbec1558-c992-4de5-91c3-4ac90e5ffec0.png���S��i���S��>�����TJA� )��:��8I)�����Ox?�������~gؙ�$���@ �����#_>z' �1���<��K������������1I�n�g����q�~�����r��q�?�g�����VS1*8($Me�^]9�{ؐ���D7-;��ݣp����ԸT%�Q���%�B�ބqT��|>Z::o��x�A�4�3:߸�(ep�t����� ô�r���7�][7��G�ч���e��Ӭ��P����?�����dޏ�+3� ��O�W���U�����{���R0��Y��,��.����/ES�X��㺐��7���ZO���qlll_I�
XZY�ɩ�������/�?�?Dof 1�͏��>5U6w8��&(�l(�K��*�iyH��MU29��=�,���N�z|��;"��sQ�\BJ�<P�����kt�S"�*��ǘN�F,#�O}�T
kO��0?��s\�#������k(��u�д�F���]:���	׹b�w�)�5��b�r���D6x���NT�n�O��r�f��a���������JR�1m����СUPJ��1�6_��]���~Z���.����B2��Ŗ�
�S���Pp$q��%�O�k��[�ph%T�v<=9M#*����[2��}qA����h�!�0TT@���IC}o����	��� \Wv��v�霾�n��G����H���ե�ہ,2�D̍�Mhq�p�A�c�.P�~�ϛ�S	��E�F�,��J�:��@�EA�=��u@&�I�5���o�sg���J	���q`\y�#t+K��7��&8&�s8��$��ag�bY����L�:)p������m��9QG n>wU��	1cYNoqc�������'9����H�o�����(�:��_y��YS'��K��($H�XJ���Ox��\0Kr�DF�>J����z�?�7E�:�0������If��'S�6����Z��j�)��qZ(�>Tѻbz�_�J�K��sX��7vF�T��:P1������vf�C�a��+��,dK)�#���@�dy�\�ͫ2��zKB���\�,����2r�<�_u��^�U*�!��6ut-w5����e	L��)i�KG��I�L�r�S���`8?E� xaaV]����0���k�\&W������s�ؽ�*�-Y��U�=Z�����[��}�xOy����:/�P���r��s��+�w��׸�b�bm�F°�(�hj�l>b�S5��)���3��Oo��/?�?]e��F�_4T�R�0�}�u���{���iѱ�2=��CS���rLm�w��TA W��5^3�>����w���bܪ����%y"Mj\�2Zim������_�$�p������~�����~�:�������׉����w3(M;�ᬣ�L�GBҗVp�i�>�V�\.���e�êJ�/-{g�>8Z�w��E��O����ȴ��N$
��b��~���z����>P��לq�И*��L���ka��BƷ�'���̰1�W�)�у��#�|~B5w�5lX� �2�߬Bo8�s���h�I���ٳ�Dՙ#��?���:�Қ��+&�6y���hk�[�f�m�b��=f�� {�q� &�
ⱊ%�Ɋ��s���3���ט#�HA,��Ӛ���"�~�8�����#���q͞2Oz�Jg��`�"��*|\R���|dÙX�z���Q�Q6|��6��𱹻�����=�baf������������w�� Ip�8WB8���9��Th��ې�<*Z��/��' ɶ��7����d��� S�//Q��O��e�O���ā>y9+UJ!E�qg��:u�����5��{�������=Ҭ�Sd�l}*V���݄����aQ\���P��jO�+���3BѰ��:Y@����a�4c���ys�x���e���{ⲳ��n�mg�n#H�c��A��`�^X+����7KTVV���(O���熇�;�6^EB�1Gtaq�0J��m/�74+���%qF�6
�>Y,���ϟS���b P��O��D���H�;/ܗ766�m�p�L�a:�u/:*,$�%#���De����L9�a�M�ۓ������DTr���������z~>�s��͘.�[L�����͏�#�	nb�,i�3���7j����j.��v���5���WB�@��f�,��,rc!�?��αuZ�w]^9F5hC�444Έ���5���32��8Y�����S�l��[Q�d�ǽ������%� ��N������s��	�����21��33��#gg�CD^|�y&ʛ��E�:�e�����T��8;�K�;I3�IF�d�-gE�ao����z
a;}{rrrXUU�ܦ(��XFN��<=\ٙ�+�\��q���pR�{#&&��������&�M��� U�lv��όD"�!� �z@A�N��Y�j���_��^yz�>I:5�3�'[1b	�3fiJ��Wb1|�J=���gs|���"VK��II�p����w`[�ۍ"n�a�'�^s6����+�-rF��H��{���u:��d?�`6�l���$��`�O-5ޣ�w�LyÚ�t�e���ί_�����0?d� �n?ɦM�;~�}�T���-.����2'�z�Z��zS����%I#Z4[)���AR��-�j���z�/x^P�|�IR�Zg�5�ҏ��S�w�����Ӻ1@�V���D�JulM�z���>2Oo%LX+�IkЏ.��,��v[��0]vv�z�{$���P��_
�j�Z ��e��D���#�ͥj�oj�z/����6�$��n��܍p��4�D:g��'/�Ϙ��h�����f��[�We�\������N�+a�^�PӸBbXE ,D��*UPV�D} ���L2e���|�L�5:�Zjim��S��F�,F�E��w�B���0�ߨ����6�K���MS��:� �5�A�__�U!H�d��q�����1�M:��b]I�svVs����2}��a�7
;��y?�7�����n���Z/�Ifz��݁��/�*,5L��@n՛�"rT�[%��Q��}MpRG�����Qj�=1�=����'!��Zm��5���������!��U�>�#�5ߥ�(3}O��[�t80� a��P������-��Pd�����Q/��>O�\V�~��v���奦�W-u��5b��Z����1�i2�s�/_�P�����1	G��ks�"r��7�%s�jYL����_K�C��ɟk:l�����Ù��sP{����B��	xkJ{E�Vn�ί�_�4Q�/���/�uY���c�����cZa,ǅY�-��W&��]����*�n��Q})뵠�-+	���ڠ� �"SS���	+�"o�o��{G�ɛ���2*+�d릑�4�Y�ɍj����?KO`�Y�
���p�I���@��߄�gb����9|��wSp�?<��=�}�:��d��S9Փh±�Y�f�2S��ͧ��0�2�ܚN~�|W�I�2��b�PU�5�~��bm�F?�	-�V�zY��.\��U�S��veZ>��L�k�����������is��^��.���yz��t圕\�H0�3A,z�:~�Z�4�5*��Z��¥�������(;c�9�V&��"�Aq�TΠ�?��,e	��i���c�-��¹��*�x!F��Y\K��1�N�!���<�ۨ፩�6��4��'����K]Q>�<熉w��V=}��O<5��.ˈ}�}���y����b���Љꉌ�rdZ��.K�4�w[񧾿vf���pq�]@�e�me���3��޲G�zCBc��6�J=�|a3Ύ��$-��`9�w	��uT�0�����QaNMm0�H�5�[��DD'��s�!�����j0�6�ͫW;��YՋ��ͳ�ɂ
���a�7r���n~:Qفs�YU@�]�������#�o�$��/�Z3by.��R*��w־s����&QU���p8<
�S]GW��7j�Miˏ�-�/�:��?��Y&���*�R�̤�v?=;��В��	�JHHX�*ڍ5*�,j-��� n7������1��l&ۿD����Y�M����F�a�L�_��=$�K�b��Չ�}�n�z���O��E�@][��)�>�J����<;;$e���3.#���Al��ǿ�0���J�;$���:j%��'5h-�v ����<0	�4z>��e�r�A)]m�k4���[p�~{}Z |'>���#L�jll���W���%73�3����L�ޫ{YJ6~u��0�L�yq�(�,���r~�|4������Pͧ!�/��#�$XC�j
����o��(A��n`�ʳ��*
���&�?���Gs4]o�t9�	��zyOH�ˋ=��×j=��Bv���&��5�߭?�:	�� �� ���k���i�L�E}Vn�Y����ϗ?��'�Vo����{X"���BM�c4��(��L鐳�@����u1#>ǧ�Lm(�a)�RXۆ4�/�~S)�
Q��	@ӱK�ISe0�pj�?��;���fS}(�p�?����O��Nl꺲�ɟ�U���֮��6C���3�p�v�i��8�����p��)k˾�Iqc���O�	R�-�dy��k���!���T�tI1�LG�*�w��)z�]y
v�\s2<*��bA�IC�.Đ�����	n�!�wd{=����ϰt�E?�<R�w�_����pE�Oa�T� ��6]$r���^������)�~e:Y�&_� ϏH�,U:��`��@-�
���Fӭ�M*m�Z�X�Ž�I�4�C���b�P�AR����.�=����5��I� zÏ�=�"�	WNt�5�z�L$��Wn@�Ḽ��K�+]�_�"Ti�_-h2�
?��(�K��0�JG׮`�H�r����bGu�#�J�TJ|Ww��8\Wj9ͨ�~,I�b
c���M�Ƒýaxh$(�6ģ�|?"�l#ļ^�w�\CڞGpV^��X�~ۯ�	��.�);v��ZZ��(��ZH}O�y��[K��>S�垎%U�!t�,�PRjg�����#�pn3����\זM�H�"w�?��&nqt8��p��)��W���L�p���up-������t��	�ęշ���$�gP;i��C��u��w�OKn�S�W:k���~�4?#S-8<2 �֟\����Ӭ��=�D�>L�W��h�����@1�PK   ���X�'k�  �  /   images/e8452abc-1b33-4025-a556-b46ce3c60df1.png��PNG

   IHDR   d   &   2r>3   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��[	�U��j{���zI��t0i�D���H$��3g<zt	G��AFe���(*3"�":.�
!,*[�$d![�ٺ�I��o����ߪ��@:�%��Mn���������zo��{r:�P$�����Jv�W��!�6Uuį��뚃�I�Op~�/���$�v�a�Pw��6�>j/��n���G�6�Tt��}l�St��~�S�J8���'����ċcÊ��h:��<���c�$�	�4@��}WM-M;0��Ј(��n�D�:��朵$��x���D����!G��t?���k�~�����]r��4�4��5��&E�NxO��i��}��\<�a&�9B�o�؈Ӹ�>�3+��ry�]T���C�ُ�ˏ@J�ìkA�e��(�϶��Έhϵ��3!��ܹ�!U�Ba�]�p!M�͜�'�Po!�8�I��sm���}瘊K��de��`?Sk�����^����i��P�"���b���LD�	��0/��ٔ��LB��:~b��*4��t����9�ae��"�K)Lȸ��t�y�GE[�e�I�Nc�W~d�⿎L}�B䉯���\a�d��V���5lL��1P]8
&]h$~�]�,��D���Wqd���t�p����1��jS�_[!b�tϣ X��B���cR�Z`�<X����2Ix��<ԧ,B�$1g�x��qV�.^��H������'N��B>�X�Dm}Y�ܰ�w�G�'f�y��h�2�r9H�	��gM��[�K_�aȧ��R�	է�fT(H��4 �^�&��P�j(Z
REx6TG�9LL1�z�RqZz4��A��"���jנ�	�W��U.P��m�ϩ��% W���ʑC�,&�� ��n#�D�j�Y��r�n����{�}�,`�@�f��I�|#̴i-T3n\>��щ�΀E�i�w$��� fϞ�k�����'.f���2A��A���~F0�'oCJ���(�Ť����j�Ѯ���h�v2�A�tt7��ۢ5I�+��>���� l^�;mC���v
%Ocڇ�N�!=z%�1���DL�����S�v���(�l�EA*�&��{;��ͨ8�MN:1t��P
�;��D� �?C�Waeft�Ǖ4�E��cČx@#f88�ȣ�&���iHU�h?�O?�$�.\H�I��4�2\��p` �H9�~�s;��/����a����0SK�*�a}V�g�F��b����&b�Al���j���A���o���	�]���VPtG�_~Ӆ�k�m���Q��`�ԃ�R��k����ކl�h���|F�5�����=�8O7����G�M����.�@�������G��Ryt&Iw؄h$	��":�%�>�Ïko��h�Q�1��H]y;ꪪn���K�޽�q0��Uo�`�RF����V�H�J�O�IT���Q�OP���$��"�
�L�k)/۵�8��6�I`ŭ�G����q8w��;y�y�������0=��D^��C��/K.,��E���4�T	�����]�<u�.���!��XJ��������7L̲ϙ�2����/���3���Y���1�"�L���%?_؞S&`�'��z�ʛl����9q,�"�d|�T	ӟ��4>��@���z�ۻ�%��!�m�w�Hr��A���+��@:�����A|���&�g����_��IÞ���u�1�y]���e�#PN"!�Q=�?��*b��;���j��i��Sf�R���F���,�aS0l��q��ڎ")(ɒ).��֧���p�Dmď�����t�CUdl>�Ep����i��5k��U��/�sd0��cv}�����m��xlk~E�wT��!̌A;�����R�o�pѠ�|-�WJ�xӨƄ�$:���H��X ym�E�R@��"����k$�:s y����1��fƺ]�8�>&^k�ϒ�G�X+�j���}�\��1�9g�^�eTo�z�`��}fnH������[qo�u���7&p��,_�4!E!�@���-˂��0MS<�w��4���4#&�>g�ْL1��]d35W"G��5̫���v�k*���֭_�K�/G�$���(b�`��T^����ά��C�;C�R�׆��Л"�9�Ag&���B��d�������4MS!Z]�444�
݋��ATWWc�̙hmmEKK��$:::��da|r��Wa�Q(`�h��Z��[�$DolCb������"�Yd�.��PY7�v*++a��0�����Khj�~�k�-|{;��e1C2��!L�

�V�x�Ј#VD0��e�SIn���V���)��kjj�`��Fz��؈T*�={���`�����*��ӧOǆ#q����c�k����y�SEL�H]&�%�m�=C͋������'��ޡ!��ރ��[a�*q�3����%��U����i��r</���l�\�.�ڱ
�)*&�E�ߧɱ:b5��:�Ţ`��g���+W
	:t������/b���طo���3Y\gFB-Y��&���M�@��*�dڞ>pS8�HӸ��B���a�����+?F�#�@	�g��N? 
&���h�˒</�k�M�;�I�ò��Ff!6Oɴ�
�^�7n��ȑ#BE]v�eصkv�܉ٳgU�u�Vq��ö�L[&~%<�� �-%�7�I"��Y��
I��
RY��W![�`���~�0�n���/aْ%�����˪��W���"����'�"�����F����Q�|j���N��Z�C���ǠdNڊ0CX-����Lٿ��f�Ē��mmm�%����=y�5Va����TY *Ո�
�j?yTgTI9�.�>2��:��[!�Ůh9��9�%��S�e-�z3�;<�� ���ݨ�6�*�Y �J���͛�x<���.tww�w�Vx��ѯ������8�3|4�O`*���0� �xW'�ɡfV�D�qp ���]��KR���6m:ló��a��������J�A��]/���"�ߎm c6��1���3��[UU%ο��jkk�!����bH$B���L{Y\�Btb�b�؅̈����	l��p2��$��E��� ��]���[��d%2��E���Q[Uq�/�o.�UV��@-_0����w�<<Sh&�0���l?]ac�c�aJd�ذ�
c;�##W�=X���0q�3���H�H*~��p�]����ds"�ۆV��ae�b [Q:k!�W}�?܃�tF��H_rl9���L���{�xte݄w�F�xU'��J�H�H8n�$�P��]��e�a/�$�y��R�2
KP]��Ϲ��zT$��y����Z�.���B!�-"g��/=$vk������G���éK9!�(/�=OpM�-��:VaO���,I�>	/�\Ċ��w�Q�Q��R��Ҕt���έ�A.o_�("���_{����}��f�~UxY%o?Čס>�?�{�~Z/���q��[��!��ea�Y�k��7L�QJd[.ֻpsh7μy����E��f(}�1¦,$r%�0�"�sk�¸�����J�w���.���_}��H]/k��4��T׌�6��؏.+�K��g����'��#��c���y�`{ ?�R�_T��X$5ў�(�.��l�Ķ�j�^�C[_��T=�����5/\��������tF}Rz��^� ������G���<E���L6V�L�퓧������;}-^'f�j�Ϛ �����EBIlPu�d�He�����8�)�𲊤�T�!�����?q�w ���#b�4�}b?$������p�|Z�P����8ht������K�N�ca���$�r�֏���<�t��,bjysJ<#��k8r�LT�,�h���y�}���Q,oCJ�_>4a{G�n [Qj�;�V�A�{�&�
U#���Zɡ\�����ק�e��gޫ�]C#�a�E���ӝi䟸��xj��` U<=b�;��7��[����f��:-���D�������8���i�i������.���7�v�rkx'��y�	xp�e=7	/��H}��I�v#u���҈؆��_T�lV�8���b/�S��i�dJ�ѕB`�;E|���t�b�e�q|Au�b�w0��f�3T��e$��׬���c΋#�s�nO������%�І^����\�d{!��Mqa�_h��u����"�4U�9�B)ً��F\r�%�'��
��kXa�&0�OQ]Hu�H.�=�c�əʹ�*���O���"����u����1(�%�"ͺ�3!�&�� ��V�~�Ex]i[��i.�[_���ދ�+V`��,�C��s0w��7�r�8O.2QC�	��/k��/�,sl���-�.X��Mq3�
�K�HNID�?�^>8(��_U����3�\9H�D��k��{�݇������-!�`(�_�����.��D�����J*k�)TV�038U���������,�����Nz۽�%�G���f�7�D��؉eq"��� ��N�6g{�,�Y#�!�Oo�}�ń�Kj��a��hy��]E#��}�uw�c�j[���_ �ę�4T�\�=uB�M8>l(5��%�&v�!�:�?�;�fy[Z�3�%�ENw�?�ݬ.80s�|���{~/G�!�a�����
Q��;q����#��A2�<�1Ln��a����,�8�p�p`J&���?��B�``�t]߲C'��v�Z�>D����ؒv�~X/ݏ�?܁���U������xO.�b��)J5ᛄ�§6>(����	o�q|�y�J��~��(8VKK���و�l,F3��S���.��	}��, ,i|�y��y��!�N�sv�z�"�N��&��k���l���a���z��#gaQ�ii� ���K�����6ࠀ�IZ!�#�l?����1��L�$�RQ��qR>>�ʛ#g�X���:1�[��&>�j��Hö�h~
2�e%&�e����P)��u�Øla���1#*�8gh&��
�wh}�P$Q��SDJݫ��d�"$	�f�CM�6(���K(�"�22�
��W@%��I�p#��C��E���-�?(#�Ȟ'ٌ����.t����)��B&<Z��:�'=~��Y��.�U�3�����!�P��yc�/�o/�]�����������I�nTV�q�G>5{�������pw׎HȤ�����>gP.V@|` ��r�	�L�0����2��~K�+R��"hOj5�U<X��dZ��O�L���:n�Bm��d�'��T�{��M铿I1�6[��`sp� f�DB�%��/#N�����a!1n!E��`��ջc=�q�}�����d��\���yMu�&�eq>kX-w2��b̟��HB�I����f��ؓ�ėV�G8R��FVF{�5�{r2"�#v�
�9��mT�H
�̔B��}ҲX�C��I�o��ICn�N8�.#k��;�2>�����6��Ǳ�`�!i˅� �]��f��q�](o��G����9�e��:Ё�S��*��b�|d��E���םX������)�؋)YT.<�<Mܻ�۽�M�W	�I�h�{�X�3��wƻ9#cS�]F|��w*�������������G������ß��go=<��c���79Gu�T�iT?�';T��G���Cf/�jJ�A&�	X������KD��'�o�
2�Iˆ��    IEND�B`�PK   ���XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   ���X��l��  S�     jsons/user_defined.json�]�r7�~�jg*�%:�_�O���7��g��RS}A�ܑI��8�Th_f�i�MJ�@@VM6��G�����_N���ɓ��Ʈ���v������'��,VK�\���W6��{�����~���e������-��ٷ//��rkX�?�7��/���^-���Օ]�|?��8O��jc�'��	eM%8fH	���F%��s�(�8��8��^/���A��Z�����Fc� V+�xCҢQH)+mͩ�KU\/p�k�:	����?���+�������]�<��d�{��\_����6�XM!�[��_�>�������[.~ܹ-�7��������ް�,���/��+�	<'���bs��߭��#'O�띛����ݻ�}���g'��a�d,��bS~#����/�
��c�"I�k��۠X6+�Ĳ��J�c�*I��c�:I�_^�K���O�FB)N�ֽ��Bi��S�i�2�/���L+����4,tL*����,,tL)����<,tL(����",t�'c��B/��K�Ş����"ibOc��iEh��YɘX���=#�s��T�a"P�i�T�a�R�i�T�a�B��Ś�T�g�D�:,u̱�j�HUa�c�Q�(U���)�;��a+C����"O��\�H�f|�L�&��J���}ƾ��k���>�B�}�]K&�f�ZpęnQ�t�b���%���C�}�^]��vqH��f?PC�s����.�(�v}F�F�e�p�ٶ� ����������툻\��b�����kk��o@w�B,�������KL<�}"��nk����.�oo�)�f�}��}�ry�>y�r?^��.�w�_λ��׫��8��-��W��z�a�}7��	���^�V?�K�.���?��2�kqV3e[�"]#R[���6�q���1̘�\KԶ��)�ղE��(�[DiSb�P�'�F")�)���us�UUt�ɭ
!:2)&�rϲ��Y$�\@A4�f��P8[��nu 4D��0���SD����J�k_햏C���T�Rm�*�cκ�.}�N[�-ˊԆZ[Tjb�İ�a�&�M�3��,6�Z����ܸ�|`���N�PU�an���r�j]�2�1�d%�F�W�R3TI&�{0̌l����� {,:J�Ͷ\o_��YD(.::�8���h�ͽ�Q�-Ν8u�����H�,ۓlde`�r����꧲S� !�ծ��-9��S.k;På�������Ǌ���%@��E�\��>�7g������d�Ӭ>,�7�+���{"��~Y����;�Խ���_�[�3�������):�ܠ�����}e׳�v��\6�aL����Lºc4��5�E�v9s�x�K^��1A���h�x���7�/����[G��ô5�%��٧��׍B��Q)��$��w	�1�{���@�������%2�q��
U�u�\5�¥s��b�@Z*YW�M�i-�r�v�DI�����C����p^.$�1Sŕ|�� �a5.D0T�\�]3-�2|D����p%}\=u��%I���ٳ������~�	2{�zvQ9sT_�٥]nF~���z�E��I�u�(�)�������Z�Qje+�]����q�%���*Qi�.B,1q�"Q��ډ��pl�u��&_�(�1L��Ά�~ �w���X�$c$(=cGd�v�Od/���=���6��mոhU���tF��.���4�XK�F����?g����Β�/'��Du��%e���X�p��Fj�
1�j~����tXJ��*TFkT�Df��*�����դlt[7��k����@I#�F�p���C�*�`}�~�^h��ےy<�YuE)��h!��<΄^�����X>�Yx��-Η�%8f�_|y�d���j���>��n���GlqO�1k*�PM���)�q�]��JZ����'�3f��8<��hD�J8����q�T
bQ+*�9<Sq9N���HZ�.*�GR��� �I��Ѭ�=��Uc�d��o
��f��~0P�B¥�/pW��Kc�u�����_6���}q�[T^��۟��PW�v!�vɶ�.��R3�;\BnE��?^"1�u��D��)]?ګ�Շ�|�˖R&�˿�D�-%"%H�H��J5�/�<���Ѷ��֩��.�w�@Sո4�E��8���_o|����+7jL~�>]������Jny풢��e����1�2ME�e���:�u"����D�i�m�c���Ma��E�,�d&�0Y��"La��E�,��?u�O��S7��s'�;���>w��j��j��j���^�tE�tE�tE�tE�tE�tE�tE�tE�tEՃ
����np��j�nv�jvW�[�/�v���٪��y�sM�iC�l²�H[ʐc��NCJ�z��S-�늷���V]��R�"+-Dm5�)�L")��PV%.��H����Zȹ��L�#�4��sr,aD��"zΥ(e�h�9�e[� T���G ��5v >l  ��ku�u H� I
͹P�¼�S위L���p<w6�`Fb���f��ZV5"UWe�T���prY[VKܴ��j*�v�w�n�]-GT�4��ia�d-��6���Jsbb�UJض2�Ne7���A-s���T��
I��k�Rr�&��\V]J�1}�f����+s2"R*���}��m?Ϲ �&�rO�:~H�> Cf�-�a +|�����m¼zs)��|!0��_]�n�ٟ��=����q��w��eӸx�Vuw:�Hd�m�P��˒���l�7��0e��]y5;�y������f���
��� ��EKY���Ԩm,F����RLQ��\�e.@,�Ɖq�⊕�� ��Y�~4u���;\Ȯ����J���EX�J�b�-�P���q�w�'�p�.'�⏝
��H�rlQq�V0���}�s�-�N>�"���䇃�q�ܪ��n��/����2�-�A��Ϋ�Ϋ�F �^m[S���x�iwt��vG��ѩ_b��E�,�d&�0Y��"La��E�,�d&�0Y��"La��E�,��Z��G`��z���3ZMٮw���;=�]n�[�ٟg�v��jv�na��{v��CQS�2ٶ�m��
Kg�{���RRLY�;��-Pj�Mm4��ϊ0d�$HXm�P�T�bJT!�b�-����չƄIR8���)K��i��2#= !$ ҶP{�X@��x�� 2g�­�@w�د��s��)L��� �(�� Rf ����( ��@���E� a5:�-J��M���D2��f��TB�hpR��=��y���ؘ������־��<L����M�S8�H�P��pqGZ��0"���V� �*��ٰ�����Yg�T����d��chr���]D8��7��-E*B��`�~�����m��@�ފS%��חo���=���Gs���q�
��MO������6ӡP�u
���/b�=�#n�0��<Lt��3�{��(�/#����J�� $���Q�=��9�@:v�k�ʁ�������97
��s���9aB�)�N��X�j�ϓ2���&�i����ć�3%Nq6�8c=H�MZF}�sbc��wQ[*B�9�1��A�t��֎��͒˦?�F�1��YJE���ۛ�T��8t=�m�@��h����{��N2Dl� nK)�ir� !�����(t}��"��CGӇt2!�)8tL}Ȉ���CGև�>!�L���!�IF�Xg�+�(qg! �=Dj�q�4�X�&��Zn�$#V(����a�Qם��[u��a�Qv�#�S{�۫9&#��z��C�(!\-@D�U���"�C���4%��!XNG�l	����3&�|���d@D����!�ʀ�Z��2"�k	d�C&��H��bW�3�" ��]�� �m/B���O��b	0{���&w�L���/qx
�g�?��c ۏe����y`�P�K��V�೽�J]�8�	6,G�s\>�&1��PL�Ў�j��0��j�ro+&%V�Wc�bM��θ�F7g�Cx�o,�1���
�<�p���,�!��D8��c�{��I"�h�����HG�9�A�nX9�p����&*��C=����#� ¡��ۛ��p�������f��9��vw��ɼ�av�1����X�0�͘�D:/x��f�n"c���6cv��f���m�=�=Yav�1�}���+u>@�/��ی��A�+��ی��A��[��m���s{j�]��H;˘�D�D�Z���02�;�҂���02�6�Ԃ��1��'�'�����4��"Lq���I�-i��О� ���2v�6��{ ��+#kc H�@�y(#�(��}�gtH�����1]�ClH���Z؀z�����mlw@��(#����IH��@#����R�C��{ ��"���<�tV����F�$��*�x�V���a<x�����a<x�����a<x��P� ���B=/C]7$�x�r���a<������㡫۽�t2�㡛ܽM��㡋ݽ}��ؗi wo+>$�x��w$ݟ�vA��� ����������OLD��.7�3@"�5�y �Ѯx�[��W��;b2@"��t��>]4�� �'@��o 3@"�hy�A2�+�x���H��w�0
��=���;�xy%yº�@p�J��wE�0J�ϧ���*F��YlYrPb_�=��5c�q>J��G�4��A������8?^�A�pj��Q�g,��B��8%c�#.h��Q249��B��8?Y�A�ph��Qrf,v<྇�����rwP�5�D���y�jJ��P˜��1c�CmsJ��G���y(�L#܇��2EJ��`݀�1c4�}���C�X}�>�G磤k2�pj��jT9(��� �}���p��PrV?�}���G������:?O��H��z�)%�.Pw����D���	9(�uZ�~��fD�\!@�����b@���͐1bP�ݰ���a@���Q��
@{o�0%F���]J�*@�������
�o���H����n2%��B��;?H�A��h��C����;?A�A�0h�������<�8���>Є�;����><��D�����8%�}��w�9(�yZ�`�qR�B|4�<'�����n0S���)���Ԏw@0}̢��&`3�@IZPg���'��'�Z� ��'�(�+�VW��T��iї|�,0|���.��GU�Ŧ	�� !$.�4��n� ��<it���GՕ���mx�f�I��T�.������ͩ)�Ҫc��������Ƙ׆�­թ�\�#%�U�F(zLe�P��AsU8�D�N�?�-�.�fm�O����$�/�]����c�R����v�q�d��a����
ڕJ�z��[��oٞ�e���-�ӝ�'ӝ��ӝ�ӝ�7�ŗgOfo>�fN�f��!}���*}ڸ\�!�Y��3
�'�[Զ�j�Ԓ����}��m#��1�P�$0��Ԉ��Dec5jL�U�ֶ6���1.5՝��#t�}b��s�2��~�j&d��G3�)<�{֡\����-�
4�c)p����_�8����O�������lW;d/K�pٶ�H뜛K�q�&��4BTB��/���:1ub��������Q��eK]�윽R�����.��b*���~~�AV�h[�M��Ѻ��7���j6�q
D�b"��/��ː���ZT[�׿Z�5v)��LSnYk'�Nd����N���?PK
   ���XR d�eu  l                  cirkitFile.jsonPK
   ���Xyɜ��  �  /             �u  images/110f4c69-ce42-4daf-8800-65b9db14e3fe.pngPK
   ���X�䓶� � /             u�  images/132fbcdf-34e4-44dc-827d-09a965026955.pngPK
   ���X��g  n  /             xF images/20eadd8b-2bcf-4996-97ef-574e0a06a30b.pngPK
   �X?Q� �h  �i  /             ,_ images/27231162-8669-47ad-b932-3d7f5563edbb.jpgPK
   ��X&�n�-u  #u  /             W� images/2a76cb7e-09fe-4529-8dba-ea35a2db28d0.pngPK
   $d�X/�iz$  �$  /             �= images/2b96fa39-ee03-40f5-a6d5-dd88ef9bf1b1.pngPK
   ��X��@� �S /             �b images/2c28e0dd-d0bf-4126-a9c2-80a014cb1784.pngPK
   ���X� ���� 
� /             �v images/38cb4f51-bc72-4d24-b782-e5d855ce8001.pngPK
   ���XMe�X&� Ú /             �- images/3a8749b6-4d34-4b13-9161-5e8eca12477c.pngPK
   $d�Xx^��6� _� /             ^� images/3c85acdc-f066-473a-bd4c-bbee71bd49cd.pngPK
   ���X�Qw�M  �M  /             �H images/4a2284cc-1baa-40d9-9462-4dabdb252300.pngPK
   ���XhT���� ċ /             ǖ images/4ee7bf8d-f382-409b-ba4b-c6cc6d91a41f.pngPK
   ���X+���  D�  /             �C images/5cebb09a-e86f-4cb2-800e-22da09d26481.pngPK
   ���X~��k�6 4 /             �� images/663b53f5-e86a-4272-a51e-f5b809259b46.pngPK
   ��X:�I��  �  /             � images/684f3f0a-9a9f-442b-bbe3-87dc70a48100.pngPK
   �X�G���j  sk  /             � images/81ad8fcd-15e9-4bfc-86b2-1d5dd79993f5.jpgPK
   ���Xd��  �   /             � images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   ���X?S��� 2� /              images/99226213-8268-43da-ade8-d9d07cfcec9f.pngPK
   ���X	��#u } /              � images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   ��X�A�x�L  �M  /             pi images/a6fbdf8e-bd4c-468a-8a96-d55269d19ee2.pngPK
   ���X$�8�l  �  /             �� images/aa130aff-16e6-4627-9689-819d55b5861f.pngPK
   ���X'�Sz�  m  /             `� images/b4b7fff7-3733-43f9-86f3-7eaab1c92eea.pngPK
   ���X$7h�!  �!  /             �� images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   ���X���]  [  /             � images/cbec1558-c992-4de5-91c3-4ac90e5ffec0.pngPK
   ���X�'k�  �  /             7 images/e8452abc-1b33-4025-a556-b46ce3c60df1.pngPK
   ���XP��/�  ǽ  /             �2 images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   ���X��l��  S�               �� jsons/user_defined.jsonPK      �	  ��   